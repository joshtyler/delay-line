--------------------------------------------------
--	TO_STDLOGIC function package
--------------------------------------------------

library	ieee;
use ieee.std_logic_1164.all;
use IEEE.Vital_Primitives.all;
use IEEE.VITAL_Timing.all;

package	std_logic_SBT is

    FUNCTION To_StdLogic       ( b : BIT               ) RETURN std_logic;
    function slv_to_integer( slv : in std_logic_vector ) return integer;
    
end std_logic_SBT;

package body std_logic_SBT is

--------------------------------------------------------------------
    FUNCTION To_StdLogic       ( b : BIT               ) RETURN std_logic IS
    BEGIN
        CASE b IS
            WHEN '0' => RETURN '0';
            WHEN '1' => RETURN '1';
        END CASE;
    END;

---------------------------------------------------------------------
    -- function to convert std_logic_vector into integer 
    function slv_to_integer (slv: in std_logic_vector ) return integer is
        variable int_val : integer;
         begin
                int_val := 0;
                for i in slv'high downto slv'low loop
                    int_val := int_val * 2;
                    if slv(i) = '1' then
                        int_val := int_val + 1;
                    end if;
                end loop;
         return int_val;
        end;
end std_logic_SBT;


--============================================================================
-- SB_CARRY 
--============================================================================


    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_unsigned.all;
    library ieee;
    use ieee.VITAL_Timing.all;
    
    
entity SB_CARRY is
Port (  I0 : in  std_logic;
        I1 : in  std_logic;
        CI : in  std_logic;
        CO : out  std_logic  );
end SB_CARRY;

architecture func of SB_CARRY is
signal CI_int :std_logic:='0';
begin
process(CI)
	begin 
	   if (CI = '1' OR CI = '0') then CI_int<=CI;
	   else CI_int<= '0';
	   end if;
  end process;

CO <= (CI_int and I0) or (CI_int and I1) or (I0 and I1);
 
end func; 


--============================================================================
-- SB_CARRY_IN_MUX 
--============================================================================

library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use IEEE.Vital_Primitives.all;
use IEEE.VITAL_Timing.all;

entity SB_CARRY_IN_MUX is
generic(C_INIT:bit_vector(1 downto 0) := "00";
--        ----------------------------------------------------------------------------------
--			--VITAL PARAMETER
--		---------------------------------------------------------------------------------
		Xon   : boolean := true;
        MsgOn : boolean := false;
        tipd_carry_init_in :VitalDelayType01:= (0.0 ns, 0.0 ns);  
        tpd_carry_init_in_carry_init_out :VitalDelayType01:= (0.0 ns, 0.0 ns));
    port ( 
	  carry_init_out  : out  std_logic;
	  carry_init_in  : in  std_logic   );
--    attribute VITAL_LEVEL0 of
--      SB_CARRY_IN_MUX : entity is true;
end SB_CARRY_IN_MUX; 
 
architecture SB_CARRY_IN_MUX_V of SB_CARRY_IN_MUX is
--  attribute VITAL_LEVEL0 of
  --  SB_CARRY_IN_MUX_V : architecture is true;
	
   signal select_bits :std_logic_vector(1 downto 0);
   signal carry_init_in_ipd : std_ulogic := 'X';
   signal carry_init_out_zd : std_ulogic := 'X';

begin
   WireDelay     : block
    begin
      VitalWireDelay (carry_init_in_ipd, carry_init_in, tipd_carry_init_in);
   end block;
---------------------------------------------------------------------------------
---- BEHAVIOR SECTION
---------------------------------------------------------------------------------	
 process(select_bits,carry_init_in_ipd)
 	begin 
 	  case select_bits is
 	     when "00"=>carry_init_out_zd<='0';
 	     when "01"=>carry_init_out_zd<='1';
 	     when "10"=>carry_init_out_zd<=carry_init_in_ipd;
--	     when "11"=>carry_init_out_zd<=carry_init_in_ipd;
	     when others =>carry_init_out_zd<='0';
	  end case;
	    
   end process;
  select_bits <= TO_STDLOGICVECTOR(C_INIT);
---------------------------------------------------------------------
----VITAL path delay
--------------------------------------------------------------------
 VITALPathDelay           : process (carry_init_in_ipd, carry_init_out_zd)
   
      variable O_GlitchData : VitalGlitchDataType;
    begin    
    VitalPathDelay01 (
      OutSignal     => carry_init_out,
      GlitchData    => O_GlitchData,
      OutSignalName => "carry_init_out",
      OutTemp       => carry_init_out_zd,
      Paths         => (0 => (carry_init_in_ipd'last_event, tpd_carry_init_in_carry_init_out, true)),
      Mode          => VitalTransport,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);
  end process; 
end SB_CARRY_IN_MUX_V; 

--============================================================================
-- SB_LUT4 
--============================================================================

    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_unsigned.all;
    
entity SB_LUT4 is
   generic(LUT_INIT:bit_vector(15 downto 0) := "1100001100111100");
   port ( 
	  O  : out  std_logic;
	  I0  : in  std_logic;
	  I1  : in  std_logic;
	  I2  : in  std_logic;
	  I3  : in  std_logic   );

end SB_LUT4; 
 
architecture func of SB_LUT4 is
signal mask :std_logic_vector(15 downto 0);
signal luts:std_logic:='0';
signal I3_in:std_logic:='0';
signal I2_in:std_logic:='0';
signal I1_in:std_logic:='0';
signal I0_in:std_logic:='0';


	function lut_mux( Cbit_in:std_logic_vector; s1:std_logic; s0:std_logic)  return std_logic is 
	variable     d: std_logic_vector(3 downto 0);       		       
	variable tmp1 : std_logic_vector(1 downto 0); 
	begin 
		d:=Cbit_in; 
		tmp1 :=TO_STDLOGICVECTOR(s1 & s0);  
		if(((s1 xor s0) = '1') or ((s1 xor s0) = '0')) then 
			case tmp1 is 
			when "00" => return d(0); 
			when "01" => return d(1); 
			when "10" => return d(2);
			when "11" => return d(3); 
			when others => return 'X'; 
			end case; 
		elsif ( (d(0) xor d(1)) = '0' and (d(2) xor d(3)) = '0' and (d(0) xor d(2)) = '0') then 
			return d(0); 
		elsif ((s1 ='0') and (d(0) = d(1))) then 
			return d(0); 
		elsif ((s1 ='1') and (d(2) = d(3))) then 
			return d(2); 	
		elsif ((s0 ='0') and (d(0) = d(2))) then 
			return d(0); 			 
		elsif ((s0 ='1') and (d(1) = d(3))) then 
			return d(1); 			 
		else 
			return 'X'; 			 	
		end if;       
	end lut_mux;

begin
 	 mask <= TO_STDLOGICVECTOR(LUT_INIT);
         O<=luts;
	 I3_in <= I3;
         I2_in <= I2;
         I1_in <= I1;
         I0_in <= I0;  

	process(I3_in,I2_in,I1_in,I0_in)
   	variable INPUTS :std_logic_vector(3 downto 0);
	variable tmp    : std_logic; 
	begin 
	       
	     tmp:=(I3_in xor I2_in xor I1_in xor I0_in); 
	     INPUTS:= TO_STDLOGICVECTOR(I3_in &  I2_in  & I1_in & I0_in);

	     if ((tmp = '0') or (tmp='1')) then 
	             case INPUTS is
		     when "0000"=>luts<= mask(0)after 0.01 ns;
		     when "0001"=>luts<= mask(1)after 0.01 ns;
		     when "0010"=>luts<= mask(2)after 0.01 ns;
		     when "0011"=>luts<= mask(3)after 0.01 ns;
		     when "0100"=>luts<= mask(4)after 0.01 ns;
		     when "0101"=>luts<= mask(5)after 0.01 ns;
		     when "0110"=>luts<= mask(6)after 0.01 ns;
		     when "0111"=>luts<= mask(7)after 0.01 ns;
		     when "1000"=>luts<= mask(8)after 0.01 ns;
		     when "1001"=>luts<= mask(9)after 0.01 ns;
		     when "1010"=>luts<= mask(10)after 0.01 ns;
		     when "1011"=>luts<= mask(11)after 0.01 ns;
		     when "1100"=>luts<= mask(12)after 0.01 ns;
		     when "1101"=>luts<= mask(13)after 0.01 ns;
		     when "1110"=>luts<= mask(14)after 0.01 ns;
		     when "1111"=>luts<= mask(15)after 0.01 ns;
		     when others=>luts<= mask(0)after 0.01 ns;
		   end case;
	     else 
		luts<= lut_mux(TO_STDLOGICVECTOR(lut_mux(mask(15 downto 12),I1_in, I0_in) & lut_mux(mask(11 downto 8),I1_in,I0_in) & lut_mux(mask(7 downto 4),I1_in,I0_in) & lut_mux(mask(3 downto 0),I1_in,I0_in)),I3_in,I2_in) ;		   		
	    end if;  	
	end process; 

end func;



--============================================================================
-- SB_DFF 
--============================================================================

    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_unsigned.all;

entity SB_DFF is
   port ( 
	  Q  : out  std_logic;
	  D  : in  std_logic;
	  C  : in  std_logic  );
	  
end SB_DFF; 
 
architecture func of SB_DFF is
  signal Q_reg : std_logic := '0';
begin
  Q <= Q_reg;
 process(C)
   begin
	  if C'event and C = '1' then
		 Q_reg <= D;
      end if;
   end process;
end  func;


--============================================================================
-- SB_DFFSR 
--============================================================================

    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_unsigned.all;

entity SB_DFFSR is
   port ( 
    R  : in  std_logic;
	  Q  : out  std_logic;
	  D  : in  std_logic;
	  C  : in  std_logic  );
	  
end SB_DFFSR; 
 
architecture func of SB_DFFSR is
  signal Q_reg : std_logic := '0';
begin
  Q <= Q_reg;
 process(C)
   begin
	  if C'event and C = '1' then
	     if R = '1'then
		        Q_reg <= '0';
		   else
		        Q_reg <= D;
       end if;
    end if;
   end process;
end  func;


--============================================================================
-- SB_DFFSS 
--============================================================================

    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_unsigned.all;

entity SB_DFFSS is
   port ( 
    S  : in  std_logic;
	  Q  : out  std_logic;
	  D  : in  std_logic;
	  C  : in  std_logic  );
	  
end SB_DFFSS; 
 
architecture func of SB_DFFSS is
  signal Q_reg : std_logic := '0';
begin
  Q <= Q_reg;
 process(C)
   begin
	  if C'event and C = '1' then
	     if S = '1'then
		        Q_reg <= '1';
		   else
		        Q_reg <= D;
       end if;
    end if;
   end process;
end  func;



--============================================================================
-- SB_DFFR 
--============================================================================

    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_unsigned.all;


entity SB_DFFR is
   port ( 
    R  : in  std_logic;
	  Q  : out  std_logic;
	  D  : in  std_logic;
	  C  : in  std_logic  );
	  
end SB_DFFR; 
 
architecture func of SB_DFFR is
  signal Q_reg : std_logic := '0';
begin
  Q <= Q_reg;
 process(C , R )
   begin
	  if (C'event and C = '1') OR (R'event and R = '1')  then
	     if R = '1'then
		        Q_reg <= '0';
		   else
		        Q_reg <= D;
       end if;
    end if;
   end process;
end  func;


--============================================================================
-- SB_DFFS 
--============================================================================

    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_unsigned.all;

entity SB_DFFS is
   port ( 
    S  : in  std_logic;
	  Q  : out  std_logic;
	  D  : in  std_logic;
	  C  : in  std_logic  );
	  
end SB_DFFS; 
 
architecture func of SB_DFFS is
  signal Q_reg : std_logic := '0';
begin
  Q <= Q_reg;
 process(C , S )
   begin
	  if (C'event and C = '1') OR (S'event and S = '1')  then
	     if S = '1'then
		        Q_reg <= '1';
		   else
		        Q_reg <= D;
       end if;
    end if;
   end process;
end  func;


--============================================================================
-- SB_DFFE 
--============================================================================

    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_unsigned.all;


entity SB_DFFE is
   port ( 
    E  : in  std_logic := 'H';
	  Q  : out  std_logic;
	  D  : in  std_logic;
	  C  : in  std_logic  );
	  
end SB_DFFE; 
 
architecture func of SB_DFFE is
  signal Q_reg : std_logic := '0';
begin
  Q <= Q_reg;
 process(C)
   begin
	  if C'event and C = '1'  then
	     if E = '1'then
		        Q_reg <= D;
		   end if;
    end if;
   end process;
end  func;


--============================================================================
-- SB_DFFESR 
--============================================================================

    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_unsigned.all;


entity SB_DFFESR is
   port ( 
    E  : in  std_logic := 'H';
    R  : in  std_logic;
	  Q  : out  std_logic;
	  D  : in  std_logic;
	  C  : in  std_logic  );
	  
end SB_DFFESR; 
 
architecture func of SB_DFFESR is
  signal Q_reg : std_logic := '0';
begin
  Q <= Q_reg;
 process(C)
   begin
	  if C'event and C = '1' then
	    if E = '1' then  
	       if R = '1'then
		          Q_reg <= '0';
		     else
		          Q_reg <= D;
       end if;
      end if;
    end if;
   end process;
end  func;


--============================================================================
-- SB_DFFESS 
--============================================================================

    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_unsigned.all;


entity SB_DFFESS is
   port ( 
    E  : in  std_logic := 'H';
    S  : in  std_logic;
	  Q  : out  std_logic;
	  D  : in  std_logic;
	  C  : in  std_logic  );
	  
end SB_DFFESS; 
 
architecture func of SB_DFFESS is
  signal Q_reg : std_logic := '0';
begin
  Q <= Q_reg;
 process(C)
   begin
	  if C'event and C = '1' then
	    if E = '1' then  
	       if S = '1'then
		          Q_reg <= '1';
		     else
		          Q_reg <= D;
       end if;
      end if;
    end if;
   end process;
end  func;


--============================================================================
-- SB_DFFER 
--============================================================================

    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_unsigned.all;


entity SB_DFFER is
   port ( 
    E  : in  std_logic := 'H';
    R  : in  std_logic;
	  Q  : out  std_logic;
	  D  : in  std_logic;
	  C  : in  std_logic  );
	  
end SB_DFFER; 
 
architecture func of SB_DFFER is
  signal Q_reg : std_logic := '0';
begin
  Q <= Q_reg;
 process(C , R )
   begin
	  if (R = '1')  then
			 Q_reg <= '0';
	  else if (C'event and C = '1') then
		if E = '1' then  
	         Q_reg <= D;
         end if;
      end if;
    end if;
   end process;
end  func;


--============================================================================
-- SB_DFFES 
--============================================================================

    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_unsigned.all;

entity SB_DFFES is
   port ( 
    E  : in  std_logic := 'H';
    S  : in  std_logic;
	  Q  : out  std_logic;
	  D  : in  std_logic;
	  C  : in  std_logic  );
	  
end SB_DFFES; 
 
architecture func of SB_DFFES is
  signal Q_reg : std_logic := '0';
begin
  Q <= Q_reg;
 process(C , S)
   begin
	  if  (S = '1')  then
	              Q_reg <= '1';
		else if (C'event and C = '1') then
			if E = '1' then
		         Q_reg <= D;
         end if;
      end if;
    end if;
   end process;
end  func;


--============================================================================
-- SB_DFFN 
--============================================================================

    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_unsigned.all;

entity SB_DFFN is
   port ( 
	  Q  : out  std_logic;
	  D  : in  std_logic;
	  C  : in  std_logic  );
	  
end SB_DFFN; 
 
architecture func of SB_DFFN is
  signal Q_reg : std_logic := '0';
begin
  Q <= Q_reg;
 process(C)
   begin
	  if C'event and C = '0' then
		 Q_reg <= D;
      end if;
   end process;
end  func;


--============================================================================
-- SB_DFFNSR 
--============================================================================

    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_unsigned.all;

entity SB_DFFNSR is
   port ( 
    R  : in  std_logic;
	  Q  : out  std_logic;
	  D  : in  std_logic;
	  C  : in  std_logic  );
	  
end SB_DFFNSR; 
 
architecture func of SB_DFFNSR is
  signal Q_reg : std_logic := '0';
begin
  Q <= Q_reg;
 process(C)
   begin
	  if C'event and C = '0' then
	     if R = '1'then
		        Q_reg <= '0';
		   else
		        Q_reg <= D;
       end if;
    end if;
   end process;
end  func;



--============================================================================
-- SB_DFFNSS 
--============================================================================

    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_unsigned.all;

	entity SB_DFFNSS is
	   port ( 
	    S  : in  std_logic;
		  Q  : out  std_logic;
		  D  : in  std_logic;
		  C  : in  std_logic  );
		  
	end SB_DFFNSS; 
	 
	architecture func of SB_DFFNSS is
	  signal Q_reg : std_logic := '0';
	begin
	  Q <= Q_reg;
	 process(C)
	   begin
		  if C'event and C = '0' then
		     if S = '1'then
			        Q_reg <= '1';
			   else
			        Q_reg <= D;
	       end if;
	    end if;
	   end process;
	end  func;
	

--============================================================================
-- SB_DFFNR 
--============================================================================

    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_unsigned.all;

entity SB_DFFNR is
   port ( 
    R  : in  std_logic;
	  Q  : out  std_logic;
	  D  : in  std_logic;
	  C  : in  std_logic  );
	  
end SB_DFFNR; 
 
architecture func of SB_DFFNR is
  signal Q_reg : std_logic := '0';
begin
  Q <= Q_reg;
 process(C , R )
   begin
	  if (C'event and C = '0') OR (R'event and R = '1')  then
	     if R = '1'then
		        Q_reg <= '0';
		   else
		        Q_reg <= D;
       end if;
    end if;
   end process;
end  func;


--============================================================================
-- SB_DFFNS 
--============================================================================

    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_unsigned.all;


entity SB_DFFNS is
   port ( 
    S  : in  std_logic;
	  Q  : out  std_logic;
	  D  : in  std_logic;
	  C  : in  std_logic  );
	  
end SB_DFFNS; 
 
architecture func of SB_DFFNS is
  signal Q_reg : std_logic := '0';
begin
  Q <= Q_reg;
 process(C , S )
   begin
	  if (C'event and C = '0') OR (S'event and S = '1')  then
	     if S = '1'then
		        Q_reg <= '1';
		   else
		        Q_reg <= D;
       end if;
    end if;
   end process;
end  func;


--============================================================================
-- SB_DFFNE 
--============================================================================

    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_unsigned.all;


entity SB_DFFNE is
   port ( 
    E  : in  std_logic := 'H';
	  Q  : out  std_logic;
	  D  : in  std_logic;
	  C  : in  std_logic  );
	  
end SB_DFFNE; 
 
architecture func of SB_DFFNE is
  signal Q_reg : std_logic := '0';
begin
  Q <= Q_reg;
 process(C)
   begin
	  if C'event and C = '0'  then
	     if E = '1'then
		        Q_reg <= D;
		   end if;
    end if;
   end process;
end  func;


--============================================================================
-- SB_DFFNESR 
--============================================================================

    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_unsigned.all;


entity SB_DFFNESR is
   port ( 
    E  : in  std_logic := 'H';
    R  : in  std_logic;
	  Q  : out  std_logic;
	  D  : in  std_logic;
	  C  : in  std_logic  );
	  
end SB_DFFNESR; 
 
architecture func of SB_DFFNESR is
  signal Q_reg : std_logic := '0';
begin
  Q <= Q_reg;
 process(C)
   begin
	  if C'event and C = '0' then
	    if E = '1' then  
	       if R = '1'then
		          Q_reg <= '0';
		     else
		          Q_reg <= D;
       end if;
      end if;
    end if;
   end process;
end  func;


--============================================================================
-- SB_DFFNESS 
--============================================================================

    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_unsigned.all;



entity SB_DFFNESS is
   port ( 
    E  : in  std_logic := 'H';
    S  : in  std_logic;
	  Q  : out  std_logic;
	  D  : in  std_logic;
	  C  : in  std_logic  );
	  
end SB_DFFNESS; 
 
architecture func of SB_DFFNESS is
  signal Q_reg : std_logic := '0';
begin
  Q <= Q_reg;
 process(C)
   begin
	  if C'event and C = '0' then
	    if E = '1' then  
	       if S = '1'then
		          Q_reg <= '1';
		     else
		          Q_reg <= D;
       end if;
      end if;
    end if;
   end process;
end  func;


--============================================================================
-- SB_DFFNER 
--============================================================================

    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_unsigned.all;


entity SB_DFFNER is
   port ( 
    E  : in  std_logic := 'H';
    R  : in  std_logic;
	  Q  : out  std_logic;
	  D  : in  std_logic;
	  C  : in  std_logic  );
	  
end SB_DFFNER; 
 
architecture func of SB_DFFNER is
  signal Q_reg : std_logic := '0';
begin
  Q <= Q_reg;
 process(C , R )
   begin
	  if (R = '1')  then
			 Q_reg <= '0';
	  else if (C'event and C = '0') then
		if E = '1' then  
	         Q_reg <= D;
         end if;
      end if;
    end if;
   end process;
end  func;


--============================================================================
-- SB_DFFNES 
--============================================================================

    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_unsigned.all;

entity SB_DFFNES is
   port ( 
    E  : in  std_logic := 'H';
    S  : in  std_logic;
	  Q  : out  std_logic;
	  D  : in  std_logic;
	  C  : in  std_logic  );
	  
end SB_DFFNES; 
 
architecture func of SB_DFFNES is
  signal Q_reg : std_logic := '0';
begin
  Q <= Q_reg;
 process(C , S)
   begin
	  if  (S = '1')  then
	              Q_reg <= '1';
		else if (C'event and C = '0') then
			if E = '1' then
		         Q_reg <= D;
         end if;
      end if;
    end if;
   end process;
end  func;




----- CELL SB_RAM4KNRNW -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
use IEEE.VITAL_Timing.all; 
USE IEEE.numeric_std.ALL;

entity SB_RAM4KNRNW is

  generic ( 
           TimingChecksOn : boolean := true;
           Xon            : boolean := false;
           MsgOn          : boolean := false;
           
           tipd_RCLKN  : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_RCLKE : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_RE    : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_RADDR : VitalDelayArrayType01(7 downto 0)  := (others => (0 ns, 0 ns));
           tipd_WCLKN  : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_WCLKE : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_WE    : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_WADDR : VitalDelayArrayType01(7 downto 0)  := (others => (0 ns, 0 ns));
           tipd_MASK  : VitalDelayArrayType01(15 downto 0)  := (others => (0 ns, 0 ns));
           tipd_WDATA : VitalDelayArrayType01(15 downto 0)  := (others => (0 ns, 0 ns));

           tpd_RCLKN_RDATA : VitalDelayArrayType01(15 downto 0) := (others => (100 ns, 100 ns));

           tsetup_RADDR_RCLKN_negedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           tsetup_RADDR_RCLKN_posedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           tsetup_RCLKE_RCLKN_negedge_posedge : VitalDelayType                   := 0 ns;
           tsetup_RCLKE_RCLKN_posedge_posedge : VitalDelayType                   := 0 ns;
           tsetup_RE_RCLKN_negedge_posedge    : VitalDelayType                   := 0 ns;
           tsetup_RE_RCLKN_posedge_posedge    : VitalDelayType                   := 0 ns;

           tsetup_WADDR_WCLKN_negedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           tsetup_WADDR_WCLKN_posedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           tsetup_WDATA_WCLKN_negedge_posedge : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           tsetup_WDATA_WCLKN_posedge_posedge : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           tsetup_WCLKE_WCLKN_negedge_posedge : VitalDelayType                   := 0 ns;
           tsetup_WCLKE_WCLKN_posedge_posedge : VitalDelayType                   := 0 ns;
           tsetup_WE_WCLKN_negedge_posedge    : VitalDelayType                   := 0 ns;
           tsetup_WE_WCLKN_posedge_posedge    : VitalDelayType                   := 0 ns;
           tsetup_MASK_WCLKN_negedge_posedge  : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           tsetup_MASK_WCLKN_posedge_posedge  : VitalDelayArrayType(15 downto 0) := (others => 0 ns);

           thold_RADDR_RCLKN_negedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           thold_RADDR_RCLKN_posedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           thold_RCLKE_RCLKN_negedge_posedge : VitalDelayType                   := 0 ns;
           thold_RCLKE_RCLKN_posedge_posedge : VitalDelayType                   := 0 ns;
           thold_RE_RCLKN_negedge_posedge    : VitalDelayType                   := 0 ns;
           thold_RE_RCLKN_posedge_posedge    : VitalDelayType                   := 0 ns;

           thold_WADDR_WCLKN_negedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           thold_WADDR_WCLKN_posedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           thold_WDATA_WCLKN_negedge_posedge : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           thold_WDATA_WCLKN_posedge_posedge : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           thold_WCLKE_WCLKN_negedge_posedge : VitalDelayType                   := 0 ns;
           thold_WCLKE_WCLKN_posedge_posedge : VitalDelayType                   := 0 ns;
           thold_WE_WCLKN_negedge_posedge    : VitalDelayType                   := 0 ns;
           thold_WE_WCLKN_posedge_posedge    : VitalDelayType                   := 0 ns;
           thold_MASK_WCLKN_negedge_posedge  : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           thold_MASK_WCLKN_posedge_posedge  : VitalDelayArrayType(15 downto 0) := (others => 0 ns);

           tpw_RCLKN_negedge : VitalDelayType := 0 ns;
           tpw_RCLKN_posedge : VitalDelayType := 0 ns;
           tpw_WCLKN_negedge : VitalDelayType := 0 ns;
           tpw_WCLKN_posedge : VitalDelayType := 0 ns;

           trecovery_RCLKN_WCLKN_posedge_posedge  : VitalDelayType                   := 0 ns;
           trecovery_RCLKN_WCLKN_negedge_posedge  : VitalDelayType                   := 0 ns;
           tremoval_RCLKN_WCLKN_posedge_posedge   : VitalDelayType                   := 0 ns;
           tremoval_RCLKN_WCLKN_negedge_posedge   : VitalDelayType                   := 0 ns;
           trecovery_WCLKN_RCLKN_posedge_posedge  : VitalDelayType                   := 0 ns;
           trecovery_WCLKN_RCLKN_negedge_posedge  : VitalDelayType                   := 0 ns;
           tremoval_WCLKN_RCLKN_posedge_posedge   : VitalDelayType                   := 0 ns;
           tremoval_WCLKN_RCLKN_negedge_posedge   : VitalDelayType                   := 0 ns;


           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 15  downto 0) ;
                RCLKN  : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'L';
                RADDR : in  std_logic_vector( 7  downto 0) ;
                WCLKN  : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'L';
                WADDR : in  std_logic_vector( 7  downto 0) ;
                MASK  : in  std_logic_vector( 15  downto 0) ;
                WDATA : in  std_logic_vector( 15  downto 0)
               );
  
  --attribute VITAL_LEVEL0 of SB_RAM4KNRNW : entity is TRUE;
  
end SB_RAM4KNRNW;



architecture SB_RAM4KNRNW_V of SB_RAM4KNRNW is
    
  --attribute VITAL_LEVEL0 of SB_RAM4KNRNW_V : architecture is TRUE;

  --signal RDATA_reg : std_logic_vector( 15  downto 0) := (others => '0');

  signal MEM : std_logic_vector(4095 downto 0) ;
  signal Address_Collision_Detected : std_logic ;


  signal RADDR_ipd : std_logic_vector(7 downto 0)  := (others => 'X');
  signal RCLKN_ipd  : std_logic                    := 'X';
  signal RCLKE_ipd : std_logic                    := 'X';
  signal RE_ipd    : std_logic                    := 'X';

  signal WADDR_ipd : std_logic_vector(7 downto 0)  := (others => 'X');
  signal WCLKN_ipd  : std_logic                    := 'X';  
  signal WCLKE_ipd : std_logic                    := 'X';
  signal WE_ipd    : std_logic                    := 'X';
  signal MASK_ipd  : std_logic_vector(15 downto 0) := (others => 'X');
  signal WDATA_ipd : std_logic_vector(15 downto 0) := (others => 'X');

  signal RADDR_in : integer range 0 to 255 ;
  signal WADDR_in : integer range 0 to 255 ;

begin

  --RDATA <= RDATA_reg;

---------------------
--  Input Wire Delay
---------------------
  WireDelay : block
  begin
    RADDR_DELAY : for i in 7 downto 0 generate
       VitalWireDelay (RADDR_ipd(i), RADDR(i), tipd_RADDR(i));
    end generate RADDR_DELAY;
    VitalWireDelay (RCLKN_ipd, RCLKN, tipd_RCLKN);
    VitalWireDelay (RCLKE_ipd, RCLKE, tipd_RCLKE);
    VitalWireDelay (RE_ipd, RE, tipd_RE);
    WADDR_DELAY : for i in 7 downto 0 generate
       VitalWireDelay (WADDR_ipd(i), WADDR(i), tipd_WADDR(i));
    end generate WADDR_DELAY;
    VitalWireDelay (WCLKN_ipd, WCLKN, tipd_WCLKN);
    VitalWireDelay (WCLKE_ipd, WCLKE, tipd_WCLKE);
    VitalWireDelay (WE_ipd, WE, tipd_WE);
    MASK_DELAY : for i in 15 downto 0 generate
       VitalWireDelay (MASK_ipd(i), MASK(i), tipd_MASK(i));
    end generate MASK_DELAY;
    WDATA_DELAY : for i in 15 downto 0 generate
       VitalWireDelay (WDATA_ipd(i), WDATA(i), tipd_WDATA(i));
    end generate WDATA_DELAY;
  end block;

  process(RE_ipd,WE_ipd,WADDR_ipd,RADDR_ipd)
      begin
          if ( (WE_ipd = '1')  and (RE_ipd = '1') and ( WADDR_ipd = RADDR_ipd) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;
          assert (not(Address_Collision_Detected = '1'))
            report "Address_Collision"
            severity warning ;         
  end process; 



  VITALReadBehavior : process(RADDR_ipd,RCLKN_ipd,RCLKE_ipd,RE_ipd)
   
       variable Tviol_RADDR0_RCLKN_posedge : std_logic := '0';
       variable Tviol_RADDR1_RCLKN_posedge : std_logic := '0';
       variable Tviol_RADDR2_RCLKN_posedge : std_logic := '0';
       variable Tviol_RADDR3_RCLKN_posedge : std_logic := '0';
       variable Tviol_RADDR4_RCLKN_posedge : std_logic := '0';
       variable Tviol_RADDR5_RCLKN_posedge : std_logic := '0';
       variable Tviol_RADDR6_RCLKN_posedge : std_logic := '0';
       variable Tviol_RADDR7_RCLKN_posedge : std_logic := '0';
       variable Tviol_RCLKE_RCLKN_posedge  : std_logic := '0';
       variable Tviol_RE_RCLKN_posedge     : std_logic := '0';

       variable Tmkr_RADDR0_RCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR1_RCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR2_RCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR3_RCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR4_RCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR5_RCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR6_RCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR7_RCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RCLKE_RCLKN_posedge  : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RE_RCLKN_posedge     : VitalTimingDataType := VitalTimingDataInit;

       variable PViol_RCLKN : std_logic := '0';

       variable PInfo_RCLKN : VitalPeriodDataType ;

       variable Tviol_WCLKN_RCLKN_posedge : std_logic := '0';
       variable Tmkr_WCLKN_RCLKN_posedge  : VitalTimingDataType := VitalTimingDataInit ;
       variable Tviol_WCLKN_RCLKN_negedge : std_logic := '0';
       variable Tmkr_WCLKN_RCLKN_negedge  : VitalTimingDataType := VitalTimingDataInit ;

       variable RDATA_GlitchData0  : VitalGlitchDataType;
       variable RDATA_GlitchData1  : VitalGlitchDataType;
       variable RDATA_GlitchData2  : VitalGlitchDataType;
       variable RDATA_GlitchData3  : VitalGlitchDataType;
       variable RDATA_GlitchData4  : VitalGlitchDataType;
       variable RDATA_GlitchData5  : VitalGlitchDataType;
       variable RDATA_GlitchData6  : VitalGlitchDataType;
       variable RDATA_GlitchData7  : VitalGlitchDataType;
       variable RDATA_GlitchData8  : VitalGlitchDataType;
       variable RDATA_GlitchData9  : VitalGlitchDataType;
       variable RDATA_GlitchData10 : VitalGlitchDataType;
       variable RDATA_GlitchData11 : VitalGlitchDataType;
       variable RDATA_GlitchData12 : VitalGlitchDataType;
       variable RDATA_GlitchData13 : VitalGlitchDataType;
       variable RDATA_GlitchData14 : VitalGlitchDataType;
       variable RDATA_GlitchData15 : VitalGlitchDataType;

       variable Violation     : std_logic  := '0';

       variable temp : std_logic_vector(15 downto 0) := (others => 'X');
       variable RDATA_zd : std_logic_vector(15 downto 0) := (others => 'X');

  begin

  -------------------------
  --  Functionality Section
  -------------------------
    RADDR_in <= conv_integer(RADDR_ipd) ;
  
    if (Violation = '1') then
       RDATA <= (others => 'X') ;
    elsif ( RCLKN_ipd'event and (RCLKN_ipd = '0') and (RCLKE_ipd = '1' or RCLKE_ipd = 'H') and (RE_ipd = '1') ) then
       for i in 0 to 15 loop
         temp(i) := MEM(16*RADDR_in + i ) ;
       end loop ;
    end if ; 

    --RDATA_reg <= temp ;
    RDATA <= temp ;


  ------------------------
  --  Timing Check Section
  ------------------------
    if (TimingChecksOn) then
      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR0_RCLKN_posedge,
        TimingData     => Tmkr_RADDR0_RCLKN_posedge,
        TestSignal     => RADDR_ipd(0),
        TestSignalName => "RADDR(0)",
        TestDelay      => 0 ns,
        RefSignal      => RCLKN_ipd,
        RefSignalName  => "RCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLKN_posedge_posedge(0),
        SetupLow       => tsetup_RADDR_RCLKN_negedge_posedge(0),
        HoldLow        => thold_RADDR_RCLKN_posedge_posedge(0),
        HoldHigh       => thold_RADDR_RCLKN_negedge_posedge(0),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR1_RCLKN_posedge,
        TimingData     => Tmkr_RADDR1_RCLKN_posedge,
        TestSignal     => RADDR_ipd(1),
        TestSignalName => "RADDR(1)",
        TestDelay      => 0 ns,
        RefSignal      => RCLKN_ipd,
        RefSignalName  => "RCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLKN_posedge_posedge(1),
        SetupLow       => tsetup_RADDR_RCLKN_negedge_posedge(1),
        HoldLow        => thold_RADDR_RCLKN_posedge_posedge(1),
        HoldHigh       => thold_RADDR_RCLKN_negedge_posedge(1),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR2_RCLKN_posedge,
        TimingData     => Tmkr_RADDR2_RCLKN_posedge,
        TestSignal     => RADDR_ipd(2),
        TestSignalName => "RADDR(2)",
        TestDelay      => 0 ns,
        RefSignal      => RCLKN_ipd,
        RefSignalName  => "RCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLKN_posedge_posedge(2),
        SetupLow       => tsetup_RADDR_RCLKN_negedge_posedge(2),
        HoldLow        => thold_RADDR_RCLKN_posedge_posedge(2),
        HoldHigh       => thold_RADDR_RCLKN_negedge_posedge(2),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR3_RCLKN_posedge,
        TimingData     => Tmkr_RADDR3_RCLKN_posedge,
        TestSignal     => RADDR_ipd(3),
        TestSignalName => "RADDR(3)",
        TestDelay      => 0 ns,
        RefSignal      => RCLKN_ipd,
        RefSignalName  => "RCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLKN_posedge_posedge(3),
        SetupLow       => tsetup_RADDR_RCLKN_negedge_posedge(3),
        HoldLow        => thold_RADDR_RCLKN_posedge_posedge(3),
        HoldHigh       => thold_RADDR_RCLKN_negedge_posedge(3),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR4_RCLKN_posedge,
        TimingData     => Tmkr_RADDR4_RCLKN_posedge,
        TestSignal     => RADDR_ipd(4),
        TestSignalName => "RADDR(4)",
        TestDelay      => 0 ns,
        RefSignal      => RCLKN_ipd,
        RefSignalName  => "RCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLKN_posedge_posedge(4),
        SetupLow       => tsetup_RADDR_RCLKN_negedge_posedge(4),
        HoldLow        => thold_RADDR_RCLKN_posedge_posedge(4),
        HoldHigh       => thold_RADDR_RCLKN_negedge_posedge(4),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR5_RCLKN_posedge,
        TimingData     => Tmkr_RADDR5_RCLKN_posedge,
        TestSignal     => RADDR_ipd(5),
        TestSignalName => "RADDR(5)",
        TestDelay      => 0 ns,
        RefSignal      => RCLKN_ipd,
        RefSignalName  => "RCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLKN_posedge_posedge(5),
        SetupLow       => tsetup_RADDR_RCLKN_negedge_posedge(5),
        HoldLow        => thold_RADDR_RCLKN_posedge_posedge(5),
        HoldHigh       => thold_RADDR_RCLKN_negedge_posedge(5),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR6_RCLKN_posedge,
        TimingData     => Tmkr_RADDR6_RCLKN_posedge,
        TestSignal     => RADDR_ipd(6),
        TestSignalName => "RADDR(6)",
        TestDelay      => 0 ns,
        RefSignal      => RCLKN_ipd,
        RefSignalName  => "RCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLKN_posedge_posedge(6),
        SetupLow       => tsetup_RADDR_RCLKN_negedge_posedge(6),
        HoldLow        => thold_RADDR_RCLKN_posedge_posedge(6),
        HoldHigh       => thold_RADDR_RCLKN_negedge_posedge(6),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR7_RCLKN_posedge,
        TimingData     => Tmkr_RADDR7_RCLKN_posedge,
        TestSignal     => RADDR_ipd(7),
        TestSignalName => "RADDR(7)",
        TestDelay      => 0 ns,
        RefSignal      => RCLKN_ipd,
        RefSignalName  => "RCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLKN_posedge_posedge(7),
        SetupLow       => tsetup_RADDR_RCLKN_negedge_posedge(7),
        HoldLow        => thold_RADDR_RCLKN_posedge_posedge(7),
        HoldHigh       => thold_RADDR_RCLKN_negedge_posedge(7),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_RCLKE_RCLKN_posedge,
        TimingData     => Tmkr_RCLKE_RCLKN_posedge,
        TestSignal     => RCLKE_ipd,
        TestSignalName => "RCLKE",
        TestDelay      => 0 ns,
        RefSignal      => RCLKN_ipd,
        RefSignalName  => "RCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RCLKE_RCLKN_posedge_posedge,
        SetupLow       => tsetup_RCLKE_RCLKN_negedge_posedge,
        HoldLow        => thold_RCLKE_RCLKN_posedge_posedge,
        HoldHigh       => thold_RCLKE_RCLKN_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_RE_RCLKN_posedge,
        TimingData     => Tmkr_RE_RCLKN_posedge,
        TestSignal     => RCLKN_ipd,
        TestSignalName => "RCLKN",
        TestDelay      => 0 ns,
        RefSignal      => RCLKN_ipd,
        RefSignalName  => "RCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RE_RCLKN_posedge_posedge,
        SetupLow       => tsetup_RE_RCLKN_negedge_posedge,
        HoldLow        => thold_RE_RCLKN_posedge_posedge,
        HoldHigh       => thold_RE_RCLKN_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
        

      VitalPeriodPulseCheck (
        Violation      => Pviol_RCLKN,
        PeriodData     => PInfo_RCLKN,
        TestSignal     => RCLKN_ipd,
        TestSignalName => "RCLKN",
        TestDelay      => 0 ns,
        Period         => 0 ns,
        PulseWidthHigh => tpw_RCLKN_posedge,
        PulseWidthLow  => tpw_RCLKN_negedge,
        CheckEnabled   => true,
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

     VitalRecoveryRemovalCheck (
       Violation               => Tviol_WCLKN_RCLKN_posedge,
       TimingData              => Tmkr_WCLKN_RCLKN_posedge,
       TestSignal              => WCLKN_ipd,
       TestSignalName          => "WCLKN",
       TestDelay               => 0 ns,
       RefSignal               => RCLKN_ipd,
       RefSignalName          => "RCLKN",
       RefDelay                => 0 ns,
       Recovery                => trecovery_WCLKN_RCLKN_negedge_posedge,
       Removal                 => tremoval_WCLKN_RCLKN_negedge_posedge,
       ActiveLow               => FALSE,
       CheckEnabled            => true,
       RefTransition           => 'R',
       HeaderMsg               => "/SB_RAM4KNRNW",
       Xon                     => Xon,
       MsgOn                   => MsgOn,
       MsgSeverity             => WARNING);

     VitalRecoveryRemovalCheck (
       Violation               => Tviol_WCLKN_RCLKN_negedge,
       TimingData              => Tmkr_WCLKN_RCLKN_negedge,
       TestSignal              => WCLKN_ipd,
       TestSignalName          => "WCLKN",
       TestDelay               => 0 ns,
       RefSignal               => RCLKN_ipd,
       RefSignalName          => "RCLKN",
       RefDelay                => 0 ns,
       Recovery                => trecovery_WCLKN_RCLKN_posedge_posedge,
       Removal                 => tremoval_WCLKN_RCLKN_posedge_posedge,
       ActiveLow               => FALSE,
       CheckEnabled            => true,
       RefTransition           => 'R',
       HeaderMsg               => "/SB_RAM4KNRNW",
       Xon                     => Xon,
       MsgOn                   => MsgOn,
       MsgSeverity             => WARNING);


    end if ;

    Violation  := Pviol_RCLKN or
                  Tviol_RADDR0_RCLKN_posedge or
                  Tviol_RADDR1_RCLKN_posedge or
                  Tviol_RADDR2_RCLKN_posedge or
                  Tviol_RADDR3_RCLKN_posedge or
                  Tviol_RADDR4_RCLKN_posedge or
                  Tviol_RADDR5_RCLKN_posedge or
                  Tviol_RADDR6_RCLKN_posedge or
                  Tviol_RADDR7_RCLKN_posedge or
                  Tviol_RCLKE_RCLKN_posedge or
                  Tviol_RE_RCLKN_posedge or
                  Tviol_WCLKN_RCLKN_posedge or
                  Tviol_WCLKN_RCLKN_negedge;

    RDATA_zd(0) := Violation xor RDATA_zd(0) ;
    RDATA_zd(1) := Violation xor RDATA_zd(1) ;
    RDATA_zd(2) := Violation xor RDATA_zd(2) ;
    RDATA_zd(3) := Violation xor RDATA_zd(3) ;
    RDATA_zd(4) := Violation xor RDATA_zd(4) ;
    RDATA_zd(5) := Violation xor RDATA_zd(5) ;
    RDATA_zd(6) := Violation xor RDATA_zd(6) ;
    RDATA_zd(7) := Violation xor RDATA_zd(7) ;
    RDATA_zd(8) := Violation xor RDATA_zd(8) ;
    RDATA_zd(9) := Violation xor RDATA_zd(9) ;
    RDATA_zd(10) := Violation xor RDATA_zd(10) ;
    RDATA_zd(11) := Violation xor RDATA_zd(11) ;
    RDATA_zd(12) := Violation xor RDATA_zd(12) ;
    RDATA_zd(13) := Violation xor RDATA_zd(13) ;
    RDATA_zd(14) := Violation xor RDATA_zd(14) ;
    RDATA_zd(15) := Violation xor RDATA_zd(15) ;
    
    
    
    
    
  ----------------------
  --  Path Delay Section
  ----------------------
    VitalPathDelay01 (
      OutSignal     => RDATA(0),
      GlitchData    => RDATA_GlitchData0,
      OutSignalName => "RDATA(0)",
      OutTemp       => RDATA_zd(0),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(0), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(1),
      GlitchData    => RDATA_GlitchData1,
      OutSignalName => "RDATA(1)",
      OutTemp       => RDATA_zd(1),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(1), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(2),
      GlitchData    => RDATA_GlitchData2,
      OutSignalName => "RDATA(2)",
      OutTemp       => RDATA_zd(2),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(2), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(3),
      GlitchData    => RDATA_GlitchData3,
      OutSignalName => "RDATA(3)",
      OutTemp       => RDATA_zd(3),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(3), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(4),
      GlitchData    => RDATA_GlitchData4,
      OutSignalName => "RDATA(4)",
      OutTemp       => RDATA_zd(4),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(4), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(5),
      GlitchData    => RDATA_GlitchData5,
      OutSignalName => "RDATA(5)",
      OutTemp       => RDATA_zd(5),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(5), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(6),
      GlitchData    => RDATA_GlitchData6,
      OutSignalName => "RDATA(6)",
      OutTemp       => RDATA_zd(6),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(6), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(7),
      GlitchData    => RDATA_GlitchData7,
      OutSignalName => "RDATA(7)",
      OutTemp       => RDATA_zd(7),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(7), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(8),
      GlitchData    => RDATA_GlitchData8,
      OutSignalName => "RDATA(8)",
      OutTemp       => RDATA_zd(8),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(8), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(9),
      GlitchData    => RDATA_GlitchData9,
      OutSignalName => "RDATA(9)",
      OutTemp       => RDATA_zd(9),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(9), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(10),
      GlitchData    => RDATA_GlitchData10,
      OutSignalName => "RDATA(10)",
      OutTemp       => RDATA_zd(10),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(10), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(11),
      GlitchData    => RDATA_GlitchData11,
      OutSignalName => "RDATA(11)",
      OutTemp       => RDATA_zd(11),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(11), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(12),
      GlitchData    => RDATA_GlitchData12,
      OutSignalName => "RDATA(12)",
      OutTemp       => RDATA_zd(12),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(12), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(13),
      GlitchData    => RDATA_GlitchData13,
      OutSignalName => "RDATA(13)",
      OutTemp       => RDATA_zd(13),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(13), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(14),
      GlitchData    => RDATA_GlitchData14,
      OutSignalName => "RDATA(14)",
      OutTemp       => RDATA_zd(14),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(14), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(15),
      GlitchData    => RDATA_GlitchData15,
      OutSignalName => "RDATA(15)",
      OutTemp       => RDATA_zd(15),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(15), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);


  end process VITALReadBehavior;


  VITALWriteBehavior : process(WADDR_ipd,WCLKN_ipd,WCLKE_ipd,WE_ipd)

       variable Tviol_WADDR0_WCLKN_posedge : std_logic := '0';
       variable Tviol_WADDR1_WCLKN_posedge : std_logic := '0';
       variable Tviol_WADDR2_WCLKN_posedge : std_logic := '0';
       variable Tviol_WADDR3_WCLKN_posedge : std_logic := '0';
       variable Tviol_WADDR4_WCLKN_posedge : std_logic := '0';
       variable Tviol_WADDR5_WCLKN_posedge : std_logic := '0';
       variable Tviol_WADDR6_WCLKN_posedge : std_logic := '0';
       variable Tviol_WADDR7_WCLKN_posedge : std_logic := '0';
       variable Tviol_WCLKE_WCLKN_posedge  : std_logic := '0';
       variable Tviol_WE_WCLKN_posedge     : std_logic := '0';
       variable Tviol_WDATA0_WCLKN_posedge : std_logic := '0';
       variable Tviol_WDATA1_WCLKN_posedge : std_logic := '0';
       variable Tviol_WDATA2_WCLKN_posedge : std_logic := '0';
       variable Tviol_WDATA3_WCLKN_posedge : std_logic := '0';
       variable Tviol_WDATA4_WCLKN_posedge : std_logic := '0';
       variable Tviol_WDATA5_WCLKN_posedge : std_logic := '0';
       variable Tviol_WDATA6_WCLKN_posedge : std_logic := '0';
       variable Tviol_WDATA7_WCLKN_posedge : std_logic := '0';
       variable Tviol_WDATA8_WCLKN_posedge : std_logic := '0';
       variable Tviol_WDATA9_WCLKN_posedge : std_logic := '0';
       variable Tviol_WDATA10_WCLKN_posedge : std_logic := '0';
       variable Tviol_WDATA11_WCLKN_posedge : std_logic := '0';
       variable Tviol_WDATA12_WCLKN_posedge : std_logic := '0';
       variable Tviol_WDATA13_WCLKN_posedge : std_logic := '0';
       variable Tviol_WDATA14_WCLKN_posedge : std_logic := '0';
       variable Tviol_WDATA15_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK0_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK1_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK2_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK3_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK4_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK5_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK6_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK7_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK8_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK9_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK10_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK11_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK12_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK13_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK14_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK15_WCLKN_posedge : std_logic := '0';


       variable Tmkr_WADDR0_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR1_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR2_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR3_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR4_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR5_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR6_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR7_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WCLKE_WCLKN_posedge  : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WE_WCLKN_posedge     : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA0_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA1_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA2_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA3_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA4_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA5_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA6_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA7_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA8_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA9_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA10_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA11_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA12_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA13_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA14_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA15_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK0_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK1_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK2_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK3_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK4_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK5_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK6_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK7_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK8_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK9_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK10_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK11_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK12_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK13_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK14_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK15_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;

       variable PViol_WCLKN : std_logic := '0';

       variable PInfo_WCLKN : VitalPeriodDataType := VitalPeriodDataInit;

       variable Tviol_RCLKN_WCLKN_posedge : std_logic := '0';
       variable Tmkr_RCLKN_WCLKN_posedge  : VitalTimingDataType := VitalTimingDataInit;
       variable Tviol_RCLKN_WCLKN_negedge : std_logic := '0';
       variable Tmkr_RCLKN_WCLKN_negedge  : VitalTimingDataType := VitalTimingDataInit;


       variable Violation     : std_logic  := '0';

       variable MEM_temp : std_logic_vector(4095 downto 0) := To_StdLogicVector(INIT_F) &
                                                              To_StdLogicVector(INIT_E) &
                                                              To_StdLogicVector(INIT_D) &
                                                              To_StdLogicVector(INIT_C) &
                                                              To_StdLogicVector(INIT_B) &
                                                              To_StdLogicVector(INIT_A) &
                                                              To_StdLogicVector(INIT_9) &
                                                              To_StdLogicVector(INIT_8) &
                                                              To_StdLogicVector(INIT_7) &
                                                              To_StdLogicVector(INIT_6) &
                                                              To_StdLogicVector(INIT_5) &
                                                              To_StdLogicVector(INIT_4) &
                                                              To_StdLogicVector(INIT_3) &
                                                              To_StdLogicVector(INIT_2) &
                                                              To_StdLogicVector(INIT_1) &
                                                              To_StdLogicVector(INIT_0);
       
  begin

    Violation  := Pviol_WCLKN or
                  Tviol_WADDR0_WCLKN_posedge or
                  Tviol_WADDR1_WCLKN_posedge or
                  Tviol_WADDR2_WCLKN_posedge or
                  Tviol_WADDR3_WCLKN_posedge or
                  Tviol_WADDR4_WCLKN_posedge or
                  Tviol_WADDR5_WCLKN_posedge or
                  Tviol_WADDR6_WCLKN_posedge or
                  Tviol_WADDR7_WCLKN_posedge or
                  Tviol_WCLKE_WCLKN_posedge or
                  Tviol_WE_WCLKN_posedge or
                  Tviol_WDATA0_WCLKN_posedge or
                  Tviol_WDATA1_WCLKN_posedge or
                  Tviol_WDATA2_WCLKN_posedge or
                  Tviol_WDATA3_WCLKN_posedge or
                  Tviol_WDATA4_WCLKN_posedge or
                  Tviol_WDATA5_WCLKN_posedge or
                  Tviol_WDATA6_WCLKN_posedge or
                  Tviol_WDATA7_WCLKN_posedge or
                  Tviol_WDATA8_WCLKN_posedge or
                  Tviol_WDATA9_WCLKN_posedge or
                  Tviol_WDATA10_WCLKN_posedge or
                  Tviol_WDATA11_WCLKN_posedge or
                  Tviol_WDATA12_WCLKN_posedge or
                  Tviol_WDATA13_WCLKN_posedge or
                  Tviol_WDATA14_WCLKN_posedge or
                  Tviol_WDATA15_WCLKN_posedge or
                  Tviol_MASK0_WCLKN_posedge or
                  Tviol_MASK1_WCLKN_posedge or
                  Tviol_MASK2_WCLKN_posedge or
                  Tviol_MASK3_WCLKN_posedge or
                  Tviol_MASK4_WCLKN_posedge or
                  Tviol_MASK5_WCLKN_posedge or
                  Tviol_MASK6_WCLKN_posedge or
                  Tviol_MASK7_WCLKN_posedge or
                  Tviol_MASK8_WCLKN_posedge or
                  Tviol_MASK9_WCLKN_posedge or
                  Tviol_MASK10_WCLKN_posedge or
                  Tviol_MASK11_WCLKN_posedge or
                  Tviol_MASK12_WCLKN_posedge or
                  Tviol_MASK13_WCLKN_posedge or
                  Tviol_MASK14_WCLKN_posedge or
                  Tviol_MASK15_WCLKN_posedge or
                  Tviol_RCLKN_WCLKN_posedge or
                  Tviol_RCLKN_WCLKN_negedge;
 
-------------------------
--  Functionality Section
-------------------------

    WADDR_in <= conv_integer(WADDR_ipd) ;
  
    if (Violation = '1') then
       MEM <= (others => 'X') ;
    elsif ( WCLKN_ipd'event and (WCLKN_ipd = '0') and (WCLKE_ipd = '1' or WCLKE_ipd = 'H') and (WE_ipd = '1') ) then
       for i in 0 to 15 loop
         if (MASK(i) = '0') then
            MEM_temp(16*WADDR_in + i ) := WDATA_ipd(i) ;
         end if ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;

------------------------
--  Timing Check Section
------------------------
    if (TimingChecksOn) then
      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR0_WCLKN_posedge,
        TimingData     => Tmkr_WADDR0_WCLKN_posedge,
        TestSignal     => WADDR_ipd(0),
        TestSignalName => "WADDR(0)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLKN_posedge_posedge(0),
        SetupLow       => tsetup_WADDR_WCLKN_negedge_posedge(0),
        HoldLow        => thold_WADDR_WCLKN_posedge_posedge(0),
        HoldHigh       => thold_WADDR_WCLKN_negedge_posedge(0),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR1_WCLKN_posedge,
        TimingData     => Tmkr_WADDR1_WCLKN_posedge,
        TestSignal     => WADDR_ipd(1),
        TestSignalName => "WADDR(1)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLKN_posedge_posedge(1),
        SetupLow       => tsetup_WADDR_WCLKN_negedge_posedge(1),
        HoldLow        => thold_WADDR_WCLKN_posedge_posedge(1),
        HoldHigh       => thold_WADDR_WCLKN_negedge_posedge(1),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR2_WCLKN_posedge,
        TimingData     => Tmkr_WADDR2_WCLKN_posedge,
        TestSignal     => WADDR_ipd(2),
        TestSignalName => "WADDR(2)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLKN_posedge_posedge(2),
        SetupLow       => tsetup_WADDR_WCLKN_negedge_posedge(2),
        HoldLow        => thold_WADDR_WCLKN_posedge_posedge(2),
        HoldHigh       => thold_WADDR_WCLKN_negedge_posedge(2),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR3_WCLKN_posedge,
        TimingData     => Tmkr_WADDR3_WCLKN_posedge,
        TestSignal     => WADDR_ipd(3),
        TestSignalName => "WADDR(3)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLKN_posedge_posedge(3),
        SetupLow       => tsetup_WADDR_WCLKN_negedge_posedge(3),
        HoldLow        => thold_WADDR_WCLKN_posedge_posedge(3),
        HoldHigh       => thold_WADDR_WCLKN_negedge_posedge(3),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR4_WCLKN_posedge,
        TimingData     => Tmkr_WADDR4_WCLKN_posedge,
        TestSignal     => WADDR_ipd(4),
        TestSignalName => "WADDR(4)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLKN_posedge_posedge(4),
        SetupLow       => tsetup_WADDR_WCLKN_negedge_posedge(4),
        HoldLow        => thold_WADDR_WCLKN_posedge_posedge(4),
        HoldHigh       => thold_WADDR_WCLKN_negedge_posedge(4),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR5_WCLKN_posedge,
        TimingData     => Tmkr_WADDR5_WCLKN_posedge,
        TestSignal     => WADDR_ipd(5),
        TestSignalName => "WADDR(5)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLKN_posedge_posedge(5),
        SetupLow       => tsetup_WADDR_WCLKN_negedge_posedge(5),
        HoldLow        => thold_WADDR_WCLKN_posedge_posedge(5),
        HoldHigh       => thold_WADDR_WCLKN_negedge_posedge(5),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR6_WCLKN_posedge,
        TimingData     => Tmkr_WADDR6_WCLKN_posedge,
        TestSignal     => WADDR_ipd(6),
        TestSignalName => "WADDR(6)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLKN_posedge_posedge(6),
        SetupLow       => tsetup_WADDR_WCLKN_negedge_posedge(6),
        HoldLow        => thold_WADDR_WCLKN_posedge_posedge(6),
        HoldHigh       => thold_WADDR_WCLKN_negedge_posedge(6),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR7_WCLKN_posedge,
        TimingData     => Tmkr_WADDR7_WCLKN_posedge,
        TestSignal     => WADDR_ipd(7),
        TestSignalName => "WADDR(7)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLKN_posedge_posedge(7),
        SetupLow       => tsetup_WADDR_WCLKN_negedge_posedge(7),
        HoldLow        => thold_WADDR_WCLKN_posedge_posedge(7),
        HoldHigh       => thold_WADDR_WCLKN_negedge_posedge(7),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WCLKE_WCLKN_posedge,
        TimingData     => Tmkr_WCLKE_WCLKN_posedge,
        TestSignal     => WCLKE_ipd,
        TestSignalName => "WCLKE",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WCLKE_WCLKN_posedge_posedge,
        SetupLow       => tsetup_WCLKE_WCLKN_negedge_posedge,
        HoldLow        => thold_WCLKE_WCLKN_posedge_posedge,
        HoldHigh       => thold_WCLKE_WCLKN_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WE_WCLKN_posedge,
        TimingData     => Tmkr_WE_WCLKN_posedge,
        TestSignal     => WCLKN_ipd,
        TestSignalName => "WCLKN",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WE_WCLKN_posedge_posedge,
        SetupLow       => tsetup_WE_WCLKN_negedge_posedge,
        HoldLow        => thold_WE_WCLKN_posedge_posedge,
        HoldHigh       => thold_WE_WCLKN_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
       VitalSetupHoldCheck (
        Violation      => Tviol_WDATA0_WCLKN_posedge,
        TimingData     => Tmkr_WDATA0_WCLKN_posedge,
        TestSignal     => WDATA_ipd(0),
        TestSignalName => "WDATA(0)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(0),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(0),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(0),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(0),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA1_WCLKN_posedge,
        TimingData     => Tmkr_WDATA1_WCLKN_posedge,
        TestSignal     => WDATA_ipd(1),
        TestSignalName => "WDATA(1)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(1),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(1),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(1),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(1),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA2_WCLKN_posedge,
        TimingData     => Tmkr_WDATA2_WCLKN_posedge,
        TestSignal     => WDATA_ipd(2),
        TestSignalName => "WDATA(2)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(2),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(2),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(2),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(2),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA3_WCLKN_posedge,
        TimingData     => Tmkr_WDATA3_WCLKN_posedge,
        TestSignal     => WDATA_ipd(3),
        TestSignalName => "WDATA(3)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(3),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(3),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(3),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(3),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA4_WCLKN_posedge,
        TimingData     => Tmkr_WDATA4_WCLKN_posedge,
        TestSignal     => WDATA_ipd(4),
        TestSignalName => "WDATA(4)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(4),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(4),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(4),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(4),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA5_WCLKN_posedge,
        TimingData     => Tmkr_WDATA5_WCLKN_posedge,
        TestSignal     => WDATA_ipd(5),
        TestSignalName => "WDATA(5)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(5),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(5),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(5),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(5),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA6_WCLKN_posedge,
        TimingData     => Tmkr_WDATA6_WCLKN_posedge,
        TestSignal     => WDATA_ipd(6),
        TestSignalName => "WDATA(6)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(6),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(6),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(6),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(6),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA7_WCLKN_posedge,
        TimingData     => Tmkr_WDATA7_WCLKN_posedge,
        TestSignal     => WDATA_ipd(7),
        TestSignalName => "WDATA(7)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(7),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(7),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(7),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(7),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

       VitalSetupHoldCheck (
        Violation      => Tviol_WDATA8_WCLKN_posedge,
        TimingData     => Tmkr_WDATA8_WCLKN_posedge,
        TestSignal     => WDATA_ipd(8),
        TestSignalName => "WDATA(8)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(8),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(8),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(8),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(8),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA9_WCLKN_posedge,
        TimingData     => Tmkr_WDATA9_WCLKN_posedge,
        TestSignal     => WDATA_ipd(9),
        TestSignalName => "WDATA(9)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(9),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(9),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(9),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(9),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA10_WCLKN_posedge,
        TimingData     => Tmkr_WDATA10_WCLKN_posedge,
        TestSignal     => WDATA_ipd(10),
        TestSignalName => "WDATA(10)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(10),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(10),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(10),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(10),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA11_WCLKN_posedge,
        TimingData     => Tmkr_WDATA11_WCLKN_posedge,
        TestSignal     => WDATA_ipd(11),
        TestSignalName => "WDATA(11)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(11),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(11),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(11),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(11),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA12_WCLKN_posedge,
        TimingData     => Tmkr_WDATA12_WCLKN_posedge,
        TestSignal     => WDATA_ipd(12),
        TestSignalName => "WDATA(12)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(12),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(12),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(12),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(12),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA13_WCLKN_posedge,
        TimingData     => Tmkr_WDATA13_WCLKN_posedge,
        TestSignal     => WDATA_ipd(13),
        TestSignalName => "WDATA(13)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(13),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(13),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(13),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(13),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA14_WCLKN_posedge,
        TimingData     => Tmkr_WDATA14_WCLKN_posedge,
        TestSignal     => WDATA_ipd(14),
        TestSignalName => "WDATA(14)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(14),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(14),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(14),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(14),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA15_WCLKN_posedge,
        TimingData     => Tmkr_WDATA15_WCLKN_posedge,
        TestSignal     => WDATA_ipd(15),
        TestSignalName => "WDATA(15)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(15),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(15),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(15),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(15),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

       VitalSetupHoldCheck (
        Violation      => Tviol_MASK0_WCLKN_posedge,
        TimingData     => Tmkr_MASK0_WCLKN_posedge,
        TestSignal     => MASK_ipd(0),
        TestSignalName => "MASK(0)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(0),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(0),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(0),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(0),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK1_WCLKN_posedge,
        TimingData     => Tmkr_MASK1_WCLKN_posedge,
        TestSignal     => MASK_ipd(1),
        TestSignalName => "MASK(1)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(1),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(1),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(1),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(1),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK2_WCLKN_posedge,
        TimingData     => Tmkr_MASK2_WCLKN_posedge,
        TestSignal     => MASK_ipd(2),
        TestSignalName => "MASK(2)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(2),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(2),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(2),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(2),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK3_WCLKN_posedge,
        TimingData     => Tmkr_MASK3_WCLKN_posedge,
        TestSignal     => MASK_ipd(3),
        TestSignalName => "MASK(3)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(3),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(3),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(3),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(3),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK4_WCLKN_posedge,
        TimingData     => Tmkr_MASK4_WCLKN_posedge,
        TestSignal     => MASK_ipd(4),
        TestSignalName => "MASK(4)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(4),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(4),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(4),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(4),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_MASK5_WCLKN_posedge,
        TimingData     => Tmkr_MASK5_WCLKN_posedge,
        TestSignal     => MASK_ipd(5),
        TestSignalName => "MASK(5)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(5),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(5),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(5),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(5),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_MASK6_WCLKN_posedge,
        TimingData     => Tmkr_MASK6_WCLKN_posedge,
        TestSignal     => MASK_ipd(6),
        TestSignalName => "MASK(6)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(6),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(6),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(6),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(6),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_MASK7_WCLKN_posedge,
        TimingData     => Tmkr_MASK7_WCLKN_posedge,
        TestSignal     => MASK_ipd(7),
        TestSignalName => "MASK(7)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(7),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(7),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(7),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(7),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

       VitalSetupHoldCheck (
        Violation      => Tviol_MASK8_WCLKN_posedge,
        TimingData     => Tmkr_MASK8_WCLKN_posedge,
        TestSignal     => MASK_ipd(8),
        TestSignalName => "MASK(8)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(8),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(8),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(8),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(8),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK9_WCLKN_posedge,
        TimingData     => Tmkr_MASK9_WCLKN_posedge,
        TestSignal     => MASK_ipd(9),
        TestSignalName => "MASK(9)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(9),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(9),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(9),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(9),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK10_WCLKN_posedge,
        TimingData     => Tmkr_MASK10_WCLKN_posedge,
        TestSignal     => MASK_ipd(10),
        TestSignalName => "MASK(10)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(10),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(10),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(10),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(10),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK11_WCLKN_posedge,
        TimingData     => Tmkr_MASK11_WCLKN_posedge,
        TestSignal     => MASK_ipd(11),
        TestSignalName => "MASK(11)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(11),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(11),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(11),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(11),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK12_WCLKN_posedge,
        TimingData     => Tmkr_MASK12_WCLKN_posedge,
        TestSignal     => MASK_ipd(12),
        TestSignalName => "MASK(12)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(12),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(12),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(12),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(12),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_MASK13_WCLKN_posedge,
        TimingData     => Tmkr_MASK13_WCLKN_posedge,
        TestSignal     => MASK_ipd(13),
        TestSignalName => "MASK(13)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(13),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(13),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(13),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(13),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_MASK14_WCLKN_posedge,
        TimingData     => Tmkr_MASK14_WCLKN_posedge,
        TestSignal     => MASK_ipd(14),
        TestSignalName => "MASK(14)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(14),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(14),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(14),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(14),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_MASK15_WCLKN_posedge,
        TimingData     => Tmkr_MASK15_WCLKN_posedge,
        TestSignal     => MASK_ipd(15),
        TestSignalName => "MASK(15)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(15),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(15),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(15),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(15),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
   

      VitalPeriodPulseCheck (
        Violation      => Pviol_WCLKN,
        PeriodData     => PInfo_WCLKN,
        TestSignal     => WCLKN_ipd,
        TestSignalName => "WCLKN",
        TestDelay      => 0 ns,
        Period         => 0 ns,
        PulseWidthHigh => tpw_WCLKN_posedge,
        PulseWidthLow  => tpw_WCLKN_negedge,
        CheckEnabled   => true,
        HeaderMsg      => "/SB_RAM4KNRNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);


     VitalRecoveryRemovalCheck (
       Violation               => Tviol_RCLKN_WCLKN_posedge,
       TimingData              => Tmkr_RCLKN_WCLKN_posedge,
       TestSignal              => RCLKN_ipd,
       TestSignalName          => "RCLKN",
       TestDelay               => 0 ns,
       RefSignal               => WCLKN_ipd,
       RefSignalName          => "WCLKN",
       RefDelay                => 0 ns,
       Recovery                => trecovery_RCLKN_WCLKN_negedge_posedge,
       Removal                 => tremoval_RCLKN_WCLKN_negedge_posedge,
       ActiveLow               => FALSE,
       CheckEnabled            => true,
       RefTransition           => 'R',
       HeaderMsg               => "/SB_RAM4KNRNW",
       Xon                     => Xon,
       MsgOn                   => MsgOn,
       MsgSeverity             => WARNING);

     VitalRecoveryRemovalCheck (
       Violation               => Tviol_RCLKN_WCLKN_negedge,
       TimingData              => Tmkr_RCLKN_WCLKN_negedge,
       TestSignal              => RCLKN_ipd,
       TestSignalName          => "RCLKN",
       TestDelay               => 0 ns,
       RefSignal               => WCLKN_ipd,
       RefSignalName          => "WCLKN",
       RefDelay                => 0 ns,
       Recovery                => trecovery_RCLKN_WCLKN_posedge_posedge,
       Removal                 => tremoval_WCLKN_RCLKN_posedge_posedge,
       ActiveLow               => FALSE,
       CheckEnabled            => true,
       RefTransition           => 'R',
       HeaderMsg               => "/SB_RAM4KNRNW",
       Xon                     => Xon,
       MsgOn                   => MsgOn,
       MsgSeverity             => WARNING);


    end if ;

  end process VITALWriteBehavior;

end SB_RAM4KNRNW_V;


----- CELL SB_RAM4KNW -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
use IEEE.VITAL_Timing.all; 
USE IEEE.numeric_std.ALL;

entity SB_RAM4KNW is

  generic ( 
           TimingChecksOn : boolean := true;
           Xon            : boolean := false;
           MsgOn          : boolean := false;
           
           tipd_RCLK  : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_RCLKE : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_RE    : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_RADDR : VitalDelayArrayType01(7 downto 0)  := (others => (0 ns, 0 ns));
           tipd_WCLKN  : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_WCLKE : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_WE    : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_WADDR : VitalDelayArrayType01(7 downto 0)  := (others => (0 ns, 0 ns));
           tipd_MASK  : VitalDelayArrayType01(15 downto 0)  := (others => (0 ns, 0 ns));
           tipd_WDATA : VitalDelayArrayType01(15 downto 0)  := (others => (0 ns, 0 ns));

           tpd_RCLK_RDATA : VitalDelayArrayType01(15 downto 0) := (others => (100 ns, 100 ns));
           tpd_RCLK_RDATA_posedge : VitalDelayArrayType01(15 downto 0) := (others => (100 ns, 100 ns));

           tsetup_RADDR_RCLK_negedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           tsetup_RADDR_RCLK_posedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           tsetup_RCLKE_RCLK_negedge_posedge : VitalDelayType                   := 0 ns;
           tsetup_RCLKE_RCLK_posedge_posedge : VitalDelayType                   := 0 ns;
           tsetup_RE_RCLK_negedge_posedge    : VitalDelayType                   := 0 ns;
           tsetup_RE_RCLK_posedge_posedge    : VitalDelayType                   := 0 ns;

           tsetup_WADDR_WCLKN_negedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           tsetup_WADDR_WCLKN_posedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           tsetup_WDATA_WCLKN_negedge_posedge : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           tsetup_WDATA_WCLKN_posedge_posedge : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           tsetup_WCLKE_WCLKN_negedge_posedge : VitalDelayType                   := 0 ns;
           tsetup_WCLKE_WCLKN_posedge_posedge : VitalDelayType                   := 0 ns;
           tsetup_WE_WCLKN_negedge_posedge    : VitalDelayType                   := 0 ns;
           tsetup_WE_WCLKN_posedge_posedge    : VitalDelayType                   := 0 ns;
           tsetup_MASK_WCLKN_negedge_posedge  : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           tsetup_MASK_WCLKN_posedge_posedge  : VitalDelayArrayType(15 downto 0) := (others => 0 ns);

           thold_RADDR_RCLK_negedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           thold_RADDR_RCLK_posedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           thold_RCLKE_RCLK_negedge_posedge : VitalDelayType                   := 0 ns;
           thold_RCLKE_RCLK_posedge_posedge : VitalDelayType                   := 0 ns;
           thold_RE_RCLK_negedge_posedge    : VitalDelayType                   := 0 ns;
           thold_RE_RCLK_posedge_posedge    : VitalDelayType                   := 0 ns;

           thold_WADDR_WCLKN_negedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           thold_WADDR_WCLKN_posedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           thold_WDATA_WCLKN_negedge_posedge : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           thold_WDATA_WCLKN_posedge_posedge : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           thold_WCLKE_WCLKN_negedge_posedge : VitalDelayType                   := 0 ns;
           thold_WCLKE_WCLKN_posedge_posedge : VitalDelayType                   := 0 ns;
           thold_WE_WCLKN_negedge_posedge    : VitalDelayType                   := 0 ns;
           thold_WE_WCLKN_posedge_posedge    : VitalDelayType                   := 0 ns;
           thold_MASK_WCLKN_negedge_posedge  : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           thold_MASK_WCLKN_posedge_posedge  : VitalDelayArrayType(15 downto 0) := (others => 0 ns);

           tpw_RCLK_negedge : VitalDelayType := 0 ns;
           tpw_RCLK_posedge : VitalDelayType := 0 ns;
           tpw_WCLKN_negedge : VitalDelayType := 0 ns;
           tpw_WCLKN_posedge : VitalDelayType := 0 ns;

           trecovery_RCLK_WCLKN_posedge_posedge  : VitalDelayType                   := 0 ns;
           trecovery_RCLK_WCLKN_negedge_posedge  : VitalDelayType                   := 0 ns;
           tremoval_RCLK_WCLKN_posedge_posedge   : VitalDelayType                   := 0 ns;
           tremoval_RCLK_WCLKN_negedge_posedge   : VitalDelayType                   := 0 ns;
           trecovery_WCLKN_RCLK_posedge_posedge  : VitalDelayType                   := 0 ns;
           trecovery_WCLKN_RCLK_negedge_posedge  : VitalDelayType                   := 0 ns;
           tremoval_WCLKN_RCLK_posedge_posedge   : VitalDelayType                   := 0 ns;
           tremoval_WCLKN_RCLK_negedge_posedge   : VitalDelayType                   := 0 ns;


           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 15  downto 0) ;
                RCLK  : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'L';
                RADDR : in  std_logic_vector( 7  downto 0) ;
                WCLKN  : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'L';
                WADDR : in  std_logic_vector( 7  downto 0) ;
                MASK  : in  std_logic_vector( 15  downto 0) ;
                WDATA : in  std_logic_vector( 15  downto 0)
               );
  
  --attribute VITAL_LEVEL0 of SB_RAM4KNW : entity is TRUE;
  
end SB_RAM4KNW;



architecture SB_RAM4KNW_V of SB_RAM4KNW is
    
  --attribute VITAL_LEVEL0 of SB_RAM4KNW_V : architecture is TRUE;

  --signal RDATA_reg : std_logic_vector( 15  downto 0) := (others => '0');

  signal MEM : std_logic_vector(4095 downto 0) ;
  signal Address_Collision_Detected : std_logic ;


  signal RADDR_ipd : std_logic_vector(7 downto 0)  := (others => '0');  
  signal RCLK_ipd  : std_logic                    := 'X';
  signal RCLKE_ipd : std_logic                    := 'X';
  signal RE_ipd    : std_logic                    := 'X';

  signal WADDR_ipd : std_logic_vector(7 downto 0)  := (others => 'X');
  signal WCLKN_ipd  : std_logic                    := 'X';  
  signal WCLKE_ipd : std_logic                    := 'X';
  signal WE_ipd    : std_logic                    := 'X';
  signal MASK_ipd  : std_logic_vector(15 downto 0) := (others => 'X');
  signal WDATA_ipd : std_logic_vector(15 downto 0) := (others => 'X');

  signal RADDR_in : integer range 0 to 255 ;
  signal WADDR_in : integer range 0 to 255 ;

begin

  --RDATA <= RDATA_reg;

---------------------
--  Input Wire Delay
---------------------
  WireDelay : block
  begin
    RADDR_DELAY : for i in 7 downto 0 generate
       VitalWireDelay (RADDR_ipd(i), RADDR(i), tipd_RADDR(i));
    end generate RADDR_DELAY;
    VitalWireDelay (RCLK_ipd, RCLK, tipd_RCLK);
    VitalWireDelay (RCLKE_ipd, RCLKE, tipd_RCLKE);
    VitalWireDelay (RE_ipd, RE, tipd_RE);
    WADDR_DELAY : for i in 7 downto 0 generate
       VitalWireDelay (WADDR_ipd(i), WADDR(i), tipd_WADDR(i));
    end generate WADDR_DELAY;
    VitalWireDelay (WCLKN_ipd, WCLKN, tipd_WCLKN);
    VitalWireDelay (WCLKE_ipd, WCLKE, tipd_WCLKE);
    VitalWireDelay (WE_ipd, WE, tipd_WE);
    MASK_DELAY : for i in 15 downto 0 generate
       VitalWireDelay (MASK_ipd(i), MASK(i), tipd_MASK(i));
    end generate MASK_DELAY;
    WDATA_DELAY : for i in 15 downto 0 generate
       VitalWireDelay (WDATA_ipd(i), WDATA(i), tipd_WDATA(i));
    end generate WDATA_DELAY;
  end block;

  process(RE_ipd,WE_ipd,WADDR_ipd,RADDR_ipd)
      begin
          if ( (WE_ipd = '1')  and (RE_ipd = '1') and ( WADDR_ipd = RADDR_ipd) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;
          assert (not(Address_Collision_Detected = '1'))
            report "Address_Collision"
            severity warning ;         
  end process; 



  VITALReadBehavior : process(RADDR_ipd,RCLK_ipd,RCLKE_ipd,RE_ipd)
   
       variable Tviol_RADDR0_RCLK_posedge : std_logic := '0';
       variable Tviol_RADDR1_RCLK_posedge : std_logic := '0';
       variable Tviol_RADDR2_RCLK_posedge : std_logic := '0';
       variable Tviol_RADDR3_RCLK_posedge : std_logic := '0';
       variable Tviol_RADDR4_RCLK_posedge : std_logic := '0';
       variable Tviol_RADDR5_RCLK_posedge : std_logic := '0';
       variable Tviol_RADDR6_RCLK_posedge : std_logic := '0';
       variable Tviol_RADDR7_RCLK_posedge : std_logic := '0';
       variable Tviol_RCLKE_RCLK_posedge  : std_logic := '0';
       variable Tviol_RE_RCLK_posedge     : std_logic := '0';

       variable Tmkr_RADDR0_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR1_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR2_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR3_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR4_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR5_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR6_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR7_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RCLKE_RCLK_posedge  : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RE_RCLK_posedge     : VitalTimingDataType := VitalTimingDataInit;

       variable PViol_RCLK : std_logic := '0';

       variable PInfo_RCLK : VitalPeriodDataType ;

       variable Tviol_WCLKN_RCLK_posedge : std_logic := '0';
       variable Tmkr_WCLKN_RCLK_posedge  : VitalTimingDataType := VitalTimingDataInit ;
       variable Tviol_WCLKN_RCLK_negedge : std_logic := '0';
       variable Tmkr_WCLKN_RCLK_negedge  : VitalTimingDataType := VitalTimingDataInit ;

       variable RDATA_GlitchData0  : VitalGlitchDataType;
       variable RDATA_GlitchData1  : VitalGlitchDataType;
       variable RDATA_GlitchData2  : VitalGlitchDataType;
       variable RDATA_GlitchData3  : VitalGlitchDataType;
       variable RDATA_GlitchData4  : VitalGlitchDataType;
       variable RDATA_GlitchData5  : VitalGlitchDataType;
       variable RDATA_GlitchData6  : VitalGlitchDataType;
       variable RDATA_GlitchData7  : VitalGlitchDataType;
       variable RDATA_GlitchData8  : VitalGlitchDataType;
       variable RDATA_GlitchData9  : VitalGlitchDataType;
       variable RDATA_GlitchData10 : VitalGlitchDataType;
       variable RDATA_GlitchData11 : VitalGlitchDataType;
       variable RDATA_GlitchData12 : VitalGlitchDataType;
       variable RDATA_GlitchData13 : VitalGlitchDataType;
       variable RDATA_GlitchData14 : VitalGlitchDataType;
       variable RDATA_GlitchData15 : VitalGlitchDataType;

       variable Violation     : std_logic  := '0';

       variable temp : std_logic_vector(15 downto 0) := (others => 'X');
       variable RDATA_zd : std_logic_vector(15 downto 0) := (others => 'X');

  begin

  -------------------------
  --  Functionality Section
  -------------------------
    RADDR_in <= conv_integer(RADDR_ipd) ;
  
    if (Violation = '1') then
       RDATA <= (others => 'X') ;
    elsif ( RCLK_ipd'event and (RCLK_ipd = '1') and (RCLKE_ipd = '1' or RCLKE_ipd = 'H') and (RE_ipd = '1') ) then
       for i in 0 to 15 loop
         temp(i) := MEM(16*RADDR_in + i ) ;
       end loop ;
    end if ; 

    --RDATA_reg <= temp ;
    RDATA <= temp ;


  ------------------------
  --  Timing Check Section
  ------------------------
    if (TimingChecksOn) then
      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR0_RCLK_posedge,
        TimingData     => Tmkr_RADDR0_RCLK_posedge,
        TestSignal     => RADDR_ipd(0),
        TestSignalName => "RADDR(0)",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(0),
        SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(0),
        HoldLow        => thold_RADDR_RCLK_posedge_posedge(0),
        HoldHigh       => thold_RADDR_RCLK_negedge_posedge(0),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR1_RCLK_posedge,
        TimingData     => Tmkr_RADDR1_RCLK_posedge,
        TestSignal     => RADDR_ipd(1),
        TestSignalName => "RADDR(1)",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(1),
        SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(1),
        HoldLow        => thold_RADDR_RCLK_posedge_posedge(1),
        HoldHigh       => thold_RADDR_RCLK_negedge_posedge(1),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR2_RCLK_posedge,
        TimingData     => Tmkr_RADDR2_RCLK_posedge,
        TestSignal     => RADDR_ipd(2),
        TestSignalName => "RADDR(2)",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(2),
        SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(2),
        HoldLow        => thold_RADDR_RCLK_posedge_posedge(2),
        HoldHigh       => thold_RADDR_RCLK_negedge_posedge(2),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR3_RCLK_posedge,
        TimingData     => Tmkr_RADDR3_RCLK_posedge,
        TestSignal     => RADDR_ipd(3),
        TestSignalName => "RADDR(3)",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(3),
        SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(3),
        HoldLow        => thold_RADDR_RCLK_posedge_posedge(3),
        HoldHigh       => thold_RADDR_RCLK_negedge_posedge(3),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR4_RCLK_posedge,
        TimingData     => Tmkr_RADDR4_RCLK_posedge,
        TestSignal     => RADDR_ipd(4),
        TestSignalName => "RADDR(4)",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(4),
        SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(4),
        HoldLow        => thold_RADDR_RCLK_posedge_posedge(4),
        HoldHigh       => thold_RADDR_RCLK_negedge_posedge(4),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR5_RCLK_posedge,
        TimingData     => Tmkr_RADDR5_RCLK_posedge,
        TestSignal     => RADDR_ipd(5),
        TestSignalName => "RADDR(5)",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(5),
        SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(5),
        HoldLow        => thold_RADDR_RCLK_posedge_posedge(5),
        HoldHigh       => thold_RADDR_RCLK_negedge_posedge(5),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR6_RCLK_posedge,
        TimingData     => Tmkr_RADDR6_RCLK_posedge,
        TestSignal     => RADDR_ipd(6),
        TestSignalName => "RADDR(6)",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(6),
        SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(6),
        HoldLow        => thold_RADDR_RCLK_posedge_posedge(6),
        HoldHigh       => thold_RADDR_RCLK_negedge_posedge(6),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR7_RCLK_posedge,
        TimingData     => Tmkr_RADDR7_RCLK_posedge,
        TestSignal     => RADDR_ipd(7),
        TestSignalName => "RADDR(7)",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(7),
        SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(7),
        HoldLow        => thold_RADDR_RCLK_posedge_posedge(7),
        HoldHigh       => thold_RADDR_RCLK_negedge_posedge(7),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_RCLKE_RCLK_posedge,
        TimingData     => Tmkr_RCLKE_RCLK_posedge,
        TestSignal     => RCLKE_ipd,
        TestSignalName => "RCLKE",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RCLKE_RCLK_posedge_posedge,
        SetupLow       => tsetup_RCLKE_RCLK_negedge_posedge,
        HoldLow        => thold_RCLKE_RCLK_posedge_posedge,
        HoldHigh       => thold_RCLKE_RCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_RE_RCLK_posedge,
        TimingData     => Tmkr_RE_RCLK_posedge,
        TestSignal     => RCLK_ipd,
        TestSignalName => "RCLK",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RE_RCLK_posedge_posedge,
        SetupLow       => tsetup_RE_RCLK_negedge_posedge,
        HoldLow        => thold_RE_RCLK_posedge_posedge,
        HoldHigh       => thold_RE_RCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
        

      VitalPeriodPulseCheck (
        Violation      => Pviol_RCLK,
        PeriodData     => PInfo_RCLK,
        TestSignal     => RCLK_ipd,
        TestSignalName => "RCLK",
        TestDelay      => 0 ns,
        Period         => 0 ns,
        PulseWidthHigh => tpw_RCLK_posedge,
        PulseWidthLow  => tpw_RCLK_negedge,
        CheckEnabled   => true,
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

     VitalRecoveryRemovalCheck (
       Violation               => Tviol_WCLKN_RCLK_posedge,
       TimingData              => Tmkr_WCLKN_RCLK_posedge,
       TestSignal              => WCLKN_ipd,
       TestSignalName          => "WCLKN",
       TestDelay               => 0 ns,
       RefSignal               => RCLK_ipd,
       RefSignalName          => "RCLK",
       RefDelay                => 0 ns,
       Recovery                => trecovery_WCLKN_RCLK_negedge_posedge,
       Removal                 => tremoval_WCLKN_RCLK_negedge_posedge,
       ActiveLow               => FALSE,
       CheckEnabled            => true,
       RefTransition           => 'R',
       HeaderMsg               => "/SB_RAM4KNW",
       Xon                     => Xon,
       MsgOn                   => MsgOn,
       MsgSeverity             => WARNING);

     VitalRecoveryRemovalCheck (
       Violation               => Tviol_WCLKN_RCLK_negedge,
       TimingData              => Tmkr_WCLKN_RCLK_negedge,
       TestSignal              => WCLKN_ipd,
       TestSignalName          => "WCLKN",
       TestDelay               => 0 ns,
       RefSignal               => RCLK_ipd,
       RefSignalName          => "RCLK",
       RefDelay                => 0 ns,
       Recovery                => trecovery_WCLKN_RCLK_posedge_posedge,
       Removal                 => tremoval_WCLKN_RCLK_posedge_posedge,
       ActiveLow               => FALSE,
       CheckEnabled            => true,
       RefTransition           => 'R',
       HeaderMsg               => "/SB_RAM4KNW",
       Xon                     => Xon,
       MsgOn                   => MsgOn,
       MsgSeverity             => WARNING);


    end if ;

    Violation  := Pviol_RCLK or
                  Tviol_RADDR0_RCLK_posedge or
                  Tviol_RADDR1_RCLK_posedge or
                  Tviol_RADDR2_RCLK_posedge or
                  Tviol_RADDR3_RCLK_posedge or
                  Tviol_RADDR4_RCLK_posedge or
                  Tviol_RADDR5_RCLK_posedge or
                  Tviol_RADDR6_RCLK_posedge or
                  Tviol_RADDR7_RCLK_posedge or
                  Tviol_RCLKE_RCLK_posedge or
                  Tviol_RE_RCLK_posedge or
                  Tviol_WCLKN_RCLK_posedge or
                  Tviol_WCLKN_RCLK_negedge;

    RDATA_zd(0) := Violation xor RDATA_zd(0) ;
    RDATA_zd(1) := Violation xor RDATA_zd(1) ;
    RDATA_zd(2) := Violation xor RDATA_zd(2) ;
    RDATA_zd(3) := Violation xor RDATA_zd(3) ;
    RDATA_zd(4) := Violation xor RDATA_zd(4) ;
    RDATA_zd(5) := Violation xor RDATA_zd(5) ;
    RDATA_zd(6) := Violation xor RDATA_zd(6) ;
    RDATA_zd(7) := Violation xor RDATA_zd(7) ;
    RDATA_zd(8) := Violation xor RDATA_zd(8) ;
    RDATA_zd(9) := Violation xor RDATA_zd(9) ;
    RDATA_zd(10) := Violation xor RDATA_zd(10) ;
    RDATA_zd(11) := Violation xor RDATA_zd(11) ;
    RDATA_zd(12) := Violation xor RDATA_zd(12) ;
    RDATA_zd(13) := Violation xor RDATA_zd(13) ;
    RDATA_zd(14) := Violation xor RDATA_zd(14) ;
    RDATA_zd(15) := Violation xor RDATA_zd(15) ;
    
    
    
    
    
  ----------------------
  --  Path Delay Section
  ----------------------
    VitalPathDelay01 (
      OutSignal     => RDATA(0),
      GlitchData    => RDATA_GlitchData0,
      OutSignalName => "RDATA(0)",
      OutTemp       => RDATA_zd(0),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(0), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(1),
      GlitchData    => RDATA_GlitchData1,
      OutSignalName => "RDATA(1)",
      OutTemp       => RDATA_zd(1),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(1), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(2),
      GlitchData    => RDATA_GlitchData2,
      OutSignalName => "RDATA(2)",
      OutTemp       => RDATA_zd(2),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(2), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(3),
      GlitchData    => RDATA_GlitchData3,
      OutSignalName => "RDATA(3)",
      OutTemp       => RDATA_zd(3),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(3), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(4),
      GlitchData    => RDATA_GlitchData4,
      OutSignalName => "RDATA(4)",
      OutTemp       => RDATA_zd(4),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(4), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(5),
      GlitchData    => RDATA_GlitchData5,
      OutSignalName => "RDATA(5)",
      OutTemp       => RDATA_zd(5),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(5), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(6),
      GlitchData    => RDATA_GlitchData6,
      OutSignalName => "RDATA(6)",
      OutTemp       => RDATA_zd(6),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(6), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(7),
      GlitchData    => RDATA_GlitchData7,
      OutSignalName => "RDATA(7)",
      OutTemp       => RDATA_zd(7),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(7), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(8),
      GlitchData    => RDATA_GlitchData8,
      OutSignalName => "RDATA(8)",
      OutTemp       => RDATA_zd(8),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(8), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(9),
      GlitchData    => RDATA_GlitchData9,
      OutSignalName => "RDATA(9)",
      OutTemp       => RDATA_zd(9),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(9), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(10),
      GlitchData    => RDATA_GlitchData10,
      OutSignalName => "RDATA(10)",
      OutTemp       => RDATA_zd(10),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(10), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(11),
      GlitchData    => RDATA_GlitchData11,
      OutSignalName => "RDATA(11)",
      OutTemp       => RDATA_zd(11),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(11), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(12),
      GlitchData    => RDATA_GlitchData12,
      OutSignalName => "RDATA(12)",
      OutTemp       => RDATA_zd(12),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(12), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(13),
      GlitchData    => RDATA_GlitchData13,
      OutSignalName => "RDATA(13)",
      OutTemp       => RDATA_zd(13),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(13), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(14),
      GlitchData    => RDATA_GlitchData14,
      OutSignalName => "RDATA(14)",
      OutTemp       => RDATA_zd(14),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(14), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(15),
      GlitchData    => RDATA_GlitchData15,
      OutSignalName => "RDATA(15)",
      OutTemp       => RDATA_zd(15),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(15), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);




  end process VITALReadBehavior;

  VITALWriteBehavior : process(WADDR_ipd,WCLKN_ipd,WCLKE_ipd,WE_ipd)

       variable Tviol_WADDR0_WCLKN_posedge : std_logic := '0';
       variable Tviol_WADDR1_WCLKN_posedge : std_logic := '0';
       variable Tviol_WADDR2_WCLKN_posedge : std_logic := '0';
       variable Tviol_WADDR3_WCLKN_posedge : std_logic := '0';
       variable Tviol_WADDR4_WCLKN_posedge : std_logic := '0';
       variable Tviol_WADDR5_WCLKN_posedge : std_logic := '0';
       variable Tviol_WADDR6_WCLKN_posedge : std_logic := '0';
       variable Tviol_WADDR7_WCLKN_posedge : std_logic := '0';
       variable Tviol_WCLKE_WCLKN_posedge  : std_logic := '0';
       variable Tviol_WE_WCLKN_posedge     : std_logic := '0';
       variable Tviol_WDATA0_WCLKN_posedge : std_logic := '0';
       variable Tviol_WDATA1_WCLKN_posedge : std_logic := '0';
       variable Tviol_WDATA2_WCLKN_posedge : std_logic := '0';
       variable Tviol_WDATA3_WCLKN_posedge : std_logic := '0';
       variable Tviol_WDATA4_WCLKN_posedge : std_logic := '0';
       variable Tviol_WDATA5_WCLKN_posedge : std_logic := '0';
       variable Tviol_WDATA6_WCLKN_posedge : std_logic := '0';
       variable Tviol_WDATA7_WCLKN_posedge : std_logic := '0';
       variable Tviol_WDATA8_WCLKN_posedge : std_logic := '0';
       variable Tviol_WDATA9_WCLKN_posedge : std_logic := '0';
       variable Tviol_WDATA10_WCLKN_posedge : std_logic := '0';
       variable Tviol_WDATA11_WCLKN_posedge : std_logic := '0';
       variable Tviol_WDATA12_WCLKN_posedge : std_logic := '0';
       variable Tviol_WDATA13_WCLKN_posedge : std_logic := '0';
       variable Tviol_WDATA14_WCLKN_posedge : std_logic := '0';
       variable Tviol_WDATA15_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK0_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK1_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK2_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK3_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK4_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK5_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK6_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK7_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK8_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK9_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK10_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK11_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK12_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK13_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK14_WCLKN_posedge : std_logic := '0';
       variable Tviol_MASK15_WCLKN_posedge : std_logic := '0';


       variable Tmkr_WADDR0_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR1_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR2_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR3_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR4_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR5_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR6_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR7_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WCLKE_WCLKN_posedge  : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WE_WCLKN_posedge     : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA0_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA1_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA2_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA3_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA4_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA5_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA6_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA7_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA8_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA9_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA10_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA11_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA12_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA13_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA14_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA15_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK0_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK1_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK2_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK3_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK4_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK5_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK6_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK7_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK8_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK9_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK10_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK11_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK12_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK13_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK14_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK15_WCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;

       variable PViol_WCLKN : std_logic := '0';

       variable PInfo_WCLKN : VitalPeriodDataType := VitalPeriodDataInit;

       variable Tviol_RCLK_WCLKN_posedge : std_logic := '0';
       variable Tmkr_RCLK_WCLKN_posedge  : VitalTimingDataType := VitalTimingDataInit;
       variable Tviol_RCLK_WCLKN_negedge : std_logic := '0';
       variable Tmkr_RCLK_WCLKN_negedge  : VitalTimingDataType := VitalTimingDataInit;


       variable Violation     : std_logic  := '0';

       variable MEM_temp : std_logic_vector(4095 downto 0) := To_StdLogicVector(INIT_F) &
                                                              To_StdLogicVector(INIT_E) &
                                                              To_StdLogicVector(INIT_D) &
                                                              To_StdLogicVector(INIT_C) &
                                                              To_StdLogicVector(INIT_B) &
                                                              To_StdLogicVector(INIT_A) &
                                                              To_StdLogicVector(INIT_9) &
                                                              To_StdLogicVector(INIT_8) &
                                                              To_StdLogicVector(INIT_7) &
                                                              To_StdLogicVector(INIT_6) &
                                                              To_StdLogicVector(INIT_5) &
                                                              To_StdLogicVector(INIT_4) &
                                                              To_StdLogicVector(INIT_3) &
                                                              To_StdLogicVector(INIT_2) &
                                                              To_StdLogicVector(INIT_1) &
                                                              To_StdLogicVector(INIT_0);
       
  begin

    Violation  := Pviol_WCLKN or
                  Tviol_WADDR0_WCLKN_posedge or
                  Tviol_WADDR1_WCLKN_posedge or
                  Tviol_WADDR2_WCLKN_posedge or
                  Tviol_WADDR3_WCLKN_posedge or
                  Tviol_WADDR4_WCLKN_posedge or
                  Tviol_WADDR5_WCLKN_posedge or
                  Tviol_WADDR6_WCLKN_posedge or
                  Tviol_WADDR7_WCLKN_posedge or
                  Tviol_WCLKE_WCLKN_posedge or
                  Tviol_WE_WCLKN_posedge or
                  Tviol_WDATA0_WCLKN_posedge or
                  Tviol_WDATA1_WCLKN_posedge or
                  Tviol_WDATA2_WCLKN_posedge or
                  Tviol_WDATA3_WCLKN_posedge or
                  Tviol_WDATA4_WCLKN_posedge or
                  Tviol_WDATA5_WCLKN_posedge or
                  Tviol_WDATA6_WCLKN_posedge or
                  Tviol_WDATA7_WCLKN_posedge or
                  Tviol_WDATA8_WCLKN_posedge or
                  Tviol_WDATA9_WCLKN_posedge or
                  Tviol_WDATA10_WCLKN_posedge or
                  Tviol_WDATA11_WCLKN_posedge or
                  Tviol_WDATA12_WCLKN_posedge or
                  Tviol_WDATA13_WCLKN_posedge or
                  Tviol_WDATA14_WCLKN_posedge or
                  Tviol_WDATA15_WCLKN_posedge or
                  Tviol_MASK0_WCLKN_posedge or
                  Tviol_MASK1_WCLKN_posedge or
                  Tviol_MASK2_WCLKN_posedge or
                  Tviol_MASK3_WCLKN_posedge or
                  Tviol_MASK4_WCLKN_posedge or
                  Tviol_MASK5_WCLKN_posedge or
                  Tviol_MASK6_WCLKN_posedge or
                  Tviol_MASK7_WCLKN_posedge or
                  Tviol_MASK8_WCLKN_posedge or
                  Tviol_MASK9_WCLKN_posedge or
                  Tviol_MASK10_WCLKN_posedge or
                  Tviol_MASK11_WCLKN_posedge or
                  Tviol_MASK12_WCLKN_posedge or
                  Tviol_MASK13_WCLKN_posedge or
                  Tviol_MASK14_WCLKN_posedge or
                  Tviol_MASK15_WCLKN_posedge or
                  Tviol_RCLK_WCLKN_posedge or
                  Tviol_RCLK_WCLKN_negedge;
 
-------------------------
--  Functionality Section
-------------------------

    WADDR_in <= conv_integer(WADDR_ipd) ;
  
    if (Violation = '1') then
       MEM <= (others => 'X') ;
    elsif ( WCLKN_ipd'event and (WCLKN_ipd = '0') and (WCLKE_ipd = '1' or WCLKE_ipd = 'H') and (WE_ipd = '1') ) then
       for i in 0 to 15 loop
         if (MASK(i) = '0') then
            MEM_temp(16*WADDR_in + i ) := WDATA_ipd(i) ;
         end if ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;

------------------------
--  Timing Check Section
------------------------
    if (TimingChecksOn) then
      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR0_WCLKN_posedge,
        TimingData     => Tmkr_WADDR0_WCLKN_posedge,
        TestSignal     => WADDR_ipd(0),
        TestSignalName => "WADDR(0)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLKN_posedge_posedge(0),
        SetupLow       => tsetup_WADDR_WCLKN_negedge_posedge(0),
        HoldLow        => thold_WADDR_WCLKN_posedge_posedge(0),
        HoldHigh       => thold_WADDR_WCLKN_negedge_posedge(0),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR1_WCLKN_posedge,
        TimingData     => Tmkr_WADDR1_WCLKN_posedge,
        TestSignal     => WADDR_ipd(1),
        TestSignalName => "WADDR(1)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLKN_posedge_posedge(1),
        SetupLow       => tsetup_WADDR_WCLKN_negedge_posedge(1),
        HoldLow        => thold_WADDR_WCLKN_posedge_posedge(1),
        HoldHigh       => thold_WADDR_WCLKN_negedge_posedge(1),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR2_WCLKN_posedge,
        TimingData     => Tmkr_WADDR2_WCLKN_posedge,
        TestSignal     => WADDR_ipd(2),
        TestSignalName => "WADDR(2)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLKN_posedge_posedge(2),
        SetupLow       => tsetup_WADDR_WCLKN_negedge_posedge(2),
        HoldLow        => thold_WADDR_WCLKN_posedge_posedge(2),
        HoldHigh       => thold_WADDR_WCLKN_negedge_posedge(2),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR3_WCLKN_posedge,
        TimingData     => Tmkr_WADDR3_WCLKN_posedge,
        TestSignal     => WADDR_ipd(3),
        TestSignalName => "WADDR(3)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLKN_posedge_posedge(3),
        SetupLow       => tsetup_WADDR_WCLKN_negedge_posedge(3),
        HoldLow        => thold_WADDR_WCLKN_posedge_posedge(3),
        HoldHigh       => thold_WADDR_WCLKN_negedge_posedge(3),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR4_WCLKN_posedge,
        TimingData     => Tmkr_WADDR4_WCLKN_posedge,
        TestSignal     => WADDR_ipd(4),
        TestSignalName => "WADDR(4)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLKN_posedge_posedge(4),
        SetupLow       => tsetup_WADDR_WCLKN_negedge_posedge(4),
        HoldLow        => thold_WADDR_WCLKN_posedge_posedge(4),
        HoldHigh       => thold_WADDR_WCLKN_negedge_posedge(4),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR5_WCLKN_posedge,
        TimingData     => Tmkr_WADDR5_WCLKN_posedge,
        TestSignal     => WADDR_ipd(5),
        TestSignalName => "WADDR(5)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLKN_posedge_posedge(5),
        SetupLow       => tsetup_WADDR_WCLKN_negedge_posedge(5),
        HoldLow        => thold_WADDR_WCLKN_posedge_posedge(5),
        HoldHigh       => thold_WADDR_WCLKN_negedge_posedge(5),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR6_WCLKN_posedge,
        TimingData     => Tmkr_WADDR6_WCLKN_posedge,
        TestSignal     => WADDR_ipd(6),
        TestSignalName => "WADDR(6)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLKN_posedge_posedge(6),
        SetupLow       => tsetup_WADDR_WCLKN_negedge_posedge(6),
        HoldLow        => thold_WADDR_WCLKN_posedge_posedge(6),
        HoldHigh       => thold_WADDR_WCLKN_negedge_posedge(6),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR7_WCLKN_posedge,
        TimingData     => Tmkr_WADDR7_WCLKN_posedge,
        TestSignal     => WADDR_ipd(7),
        TestSignalName => "WADDR(7)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLKN_posedge_posedge(7),
        SetupLow       => tsetup_WADDR_WCLKN_negedge_posedge(7),
        HoldLow        => thold_WADDR_WCLKN_posedge_posedge(7),
        HoldHigh       => thold_WADDR_WCLKN_negedge_posedge(7),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WCLKE_WCLKN_posedge,
        TimingData     => Tmkr_WCLKE_WCLKN_posedge,
        TestSignal     => WCLKE_ipd,
        TestSignalName => "WCLKE",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WCLKE_WCLKN_posedge_posedge,
        SetupLow       => tsetup_WCLKE_WCLKN_negedge_posedge,
        HoldLow        => thold_WCLKE_WCLKN_posedge_posedge,
        HoldHigh       => thold_WCLKE_WCLKN_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WE_WCLKN_posedge,
        TimingData     => Tmkr_WE_WCLKN_posedge,
        TestSignal     => WCLKN_ipd,
        TestSignalName => "WCLKN",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WE_WCLKN_posedge_posedge,
        SetupLow       => tsetup_WE_WCLKN_negedge_posedge,
        HoldLow        => thold_WE_WCLKN_posedge_posedge,
        HoldHigh       => thold_WE_WCLKN_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
       VitalSetupHoldCheck (
        Violation      => Tviol_WDATA0_WCLKN_posedge,
        TimingData     => Tmkr_WDATA0_WCLKN_posedge,
        TestSignal     => WDATA_ipd(0),
        TestSignalName => "WDATA(0)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(0),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(0),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(0),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(0),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA1_WCLKN_posedge,
        TimingData     => Tmkr_WDATA1_WCLKN_posedge,
        TestSignal     => WDATA_ipd(1),
        TestSignalName => "WDATA(1)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(1),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(1),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(1),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(1),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA2_WCLKN_posedge,
        TimingData     => Tmkr_WDATA2_WCLKN_posedge,
        TestSignal     => WDATA_ipd(2),
        TestSignalName => "WDATA(2)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(2),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(2),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(2),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(2),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA3_WCLKN_posedge,
        TimingData     => Tmkr_WDATA3_WCLKN_posedge,
        TestSignal     => WDATA_ipd(3),
        TestSignalName => "WDATA(3)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(3),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(3),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(3),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(3),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA4_WCLKN_posedge,
        TimingData     => Tmkr_WDATA4_WCLKN_posedge,
        TestSignal     => WDATA_ipd(4),
        TestSignalName => "WDATA(4)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(4),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(4),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(4),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(4),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA5_WCLKN_posedge,
        TimingData     => Tmkr_WDATA5_WCLKN_posedge,
        TestSignal     => WDATA_ipd(5),
        TestSignalName => "WDATA(5)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(5),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(5),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(5),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(5),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA6_WCLKN_posedge,
        TimingData     => Tmkr_WDATA6_WCLKN_posedge,
        TestSignal     => WDATA_ipd(6),
        TestSignalName => "WDATA(6)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(6),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(6),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(6),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(6),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA7_WCLKN_posedge,
        TimingData     => Tmkr_WDATA7_WCLKN_posedge,
        TestSignal     => WDATA_ipd(7),
        TestSignalName => "WDATA(7)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(7),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(7),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(7),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(7),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

       VitalSetupHoldCheck (
        Violation      => Tviol_WDATA8_WCLKN_posedge,
        TimingData     => Tmkr_WDATA8_WCLKN_posedge,
        TestSignal     => WDATA_ipd(8),
        TestSignalName => "WDATA(8)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(8),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(8),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(8),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(8),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA9_WCLKN_posedge,
        TimingData     => Tmkr_WDATA9_WCLKN_posedge,
        TestSignal     => WDATA_ipd(9),
        TestSignalName => "WDATA(9)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(9),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(9),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(9),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(9),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA10_WCLKN_posedge,
        TimingData     => Tmkr_WDATA10_WCLKN_posedge,
        TestSignal     => WDATA_ipd(10),
        TestSignalName => "WDATA(10)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(10),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(10),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(10),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(10),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA11_WCLKN_posedge,
        TimingData     => Tmkr_WDATA11_WCLKN_posedge,
        TestSignal     => WDATA_ipd(11),
        TestSignalName => "WDATA(11)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(11),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(11),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(11),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(11),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA12_WCLKN_posedge,
        TimingData     => Tmkr_WDATA12_WCLKN_posedge,
        TestSignal     => WDATA_ipd(12),
        TestSignalName => "WDATA(12)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(12),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(12),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(12),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(12),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA13_WCLKN_posedge,
        TimingData     => Tmkr_WDATA13_WCLKN_posedge,
        TestSignal     => WDATA_ipd(13),
        TestSignalName => "WDATA(13)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(13),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(13),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(13),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(13),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA14_WCLKN_posedge,
        TimingData     => Tmkr_WDATA14_WCLKN_posedge,
        TestSignal     => WDATA_ipd(14),
        TestSignalName => "WDATA(14)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(14),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(14),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(14),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(14),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA15_WCLKN_posedge,
        TimingData     => Tmkr_WDATA15_WCLKN_posedge,
        TestSignal     => WDATA_ipd(15),
        TestSignalName => "WDATA(15)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLKN_posedge_posedge(15),
        SetupLow       => tsetup_WDATA_WCLKN_negedge_posedge(15),
        HoldLow        => thold_WDATA_WCLKN_posedge_posedge(15),
        HoldHigh       => thold_WDATA_WCLKN_negedge_posedge(15),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

       VitalSetupHoldCheck (
        Violation      => Tviol_MASK0_WCLKN_posedge,
        TimingData     => Tmkr_MASK0_WCLKN_posedge,
        TestSignal     => MASK_ipd(0),
        TestSignalName => "MASK(0)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(0),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(0),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(0),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(0),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK1_WCLKN_posedge,
        TimingData     => Tmkr_MASK1_WCLKN_posedge,
        TestSignal     => MASK_ipd(1),
        TestSignalName => "MASK(1)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(1),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(1),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(1),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(1),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK2_WCLKN_posedge,
        TimingData     => Tmkr_MASK2_WCLKN_posedge,
        TestSignal     => MASK_ipd(2),
        TestSignalName => "MASK(2)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(2),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(2),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(2),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(2),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK3_WCLKN_posedge,
        TimingData     => Tmkr_MASK3_WCLKN_posedge,
        TestSignal     => MASK_ipd(3),
        TestSignalName => "MASK(3)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(3),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(3),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(3),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(3),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK4_WCLKN_posedge,
        TimingData     => Tmkr_MASK4_WCLKN_posedge,
        TestSignal     => MASK_ipd(4),
        TestSignalName => "MASK(4)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(4),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(4),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(4),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(4),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_MASK5_WCLKN_posedge,
        TimingData     => Tmkr_MASK5_WCLKN_posedge,
        TestSignal     => MASK_ipd(5),
        TestSignalName => "MASK(5)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(5),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(5),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(5),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(5),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_MASK6_WCLKN_posedge,
        TimingData     => Tmkr_MASK6_WCLKN_posedge,
        TestSignal     => MASK_ipd(6),
        TestSignalName => "MASK(6)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(6),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(6),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(6),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(6),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_MASK7_WCLKN_posedge,
        TimingData     => Tmkr_MASK7_WCLKN_posedge,
        TestSignal     => MASK_ipd(7),
        TestSignalName => "MASK(7)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(7),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(7),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(7),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(7),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

       VitalSetupHoldCheck (
        Violation      => Tviol_MASK8_WCLKN_posedge,
        TimingData     => Tmkr_MASK8_WCLKN_posedge,
        TestSignal     => MASK_ipd(8),
        TestSignalName => "MASK(8)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(8),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(8),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(8),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(8),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK9_WCLKN_posedge,
        TimingData     => Tmkr_MASK9_WCLKN_posedge,
        TestSignal     => MASK_ipd(9),
        TestSignalName => "MASK(9)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(9),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(9),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(9),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(9),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK10_WCLKN_posedge,
        TimingData     => Tmkr_MASK10_WCLKN_posedge,
        TestSignal     => MASK_ipd(10),
        TestSignalName => "MASK(10)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(10),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(10),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(10),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(10),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK11_WCLKN_posedge,
        TimingData     => Tmkr_MASK11_WCLKN_posedge,
        TestSignal     => MASK_ipd(11),
        TestSignalName => "MASK(11)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(11),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(11),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(11),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(11),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK12_WCLKN_posedge,
        TimingData     => Tmkr_MASK12_WCLKN_posedge,
        TestSignal     => MASK_ipd(12),
        TestSignalName => "MASK(12)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(12),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(12),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(12),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(12),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_MASK13_WCLKN_posedge,
        TimingData     => Tmkr_MASK13_WCLKN_posedge,
        TestSignal     => MASK_ipd(13),
        TestSignalName => "MASK(13)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(13),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(13),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(13),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(13),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_MASK14_WCLKN_posedge,
        TimingData     => Tmkr_MASK14_WCLKN_posedge,
        TestSignal     => MASK_ipd(14),
        TestSignalName => "MASK(14)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(14),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(14),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(14),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(14),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_MASK15_WCLKN_posedge,
        TimingData     => Tmkr_MASK15_WCLKN_posedge,
        TestSignal     => MASK_ipd(15),
        TestSignalName => "MASK(15)",
        TestDelay      => 0 ns,
        RefSignal      => WCLKN_ipd,
        RefSignalName  => "WCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLKN_posedge_posedge(15),
        SetupLow       => tsetup_MASK_WCLKN_negedge_posedge(15),
        HoldLow        => thold_MASK_WCLKN_posedge_posedge(15),
        HoldHigh       => thold_MASK_WCLKN_negedge_posedge(15),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
   

      VitalPeriodPulseCheck (
        Violation      => Pviol_WCLKN,
        PeriodData     => PInfo_WCLKN,
        TestSignal     => WCLKN_ipd,
        TestSignalName => "WCLKN",
        TestDelay      => 0 ns,
        Period         => 0 ns,
        PulseWidthHigh => tpw_WCLKN_posedge,
        PulseWidthLow  => tpw_WCLKN_negedge,
        CheckEnabled   => true,
        HeaderMsg      => "/SB_RAM4KNW",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);


     VitalRecoveryRemovalCheck (
       Violation               => Tviol_RCLK_WCLKN_posedge,
       TimingData              => Tmkr_RCLK_WCLKN_posedge,
       TestSignal              => RCLK_ipd,
       TestSignalName          => "RCLK",
       TestDelay               => 0 ns,
       RefSignal               => WCLKN_ipd,
       RefSignalName          => "WCLKN",
       RefDelay                => 0 ns,
       Recovery                => trecovery_RCLK_WCLKN_negedge_posedge,
       Removal                 => tremoval_RCLK_WCLKN_negedge_posedge,
       ActiveLow               => FALSE,
       CheckEnabled            => true,
       RefTransition           => 'R',
       HeaderMsg               => "/SB_RAM4KNW",
       Xon                     => Xon,
       MsgOn                   => MsgOn,
       MsgSeverity             => WARNING);

     VitalRecoveryRemovalCheck (
       Violation               => Tviol_RCLK_WCLKN_negedge,
       TimingData              => Tmkr_RCLK_WCLKN_negedge,
       TestSignal              => RCLK_ipd,
       TestSignalName          => "RCLK",
       TestDelay               => 0 ns,
       RefSignal               => WCLKN_ipd,
       RefSignalName          => "WCLKN",
       RefDelay                => 0 ns,
       Recovery                => trecovery_RCLK_WCLKN_posedge_posedge,
       Removal                 => tremoval_WCLKN_RCLK_posedge_posedge,
       ActiveLow               => FALSE,
       CheckEnabled            => true,
       RefTransition           => 'R',
       HeaderMsg               => "/SB_RAM4KNW",
       Xon                     => Xon,
       MsgOn                   => MsgOn,
       MsgSeverity             => WARNING);


    end if ;



  end process VITALWriteBehavior;



end SB_RAM4KNW_V;



----- CELL SB_RAM4KNR -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
use IEEE.VITAL_Timing.all; 
USE IEEE.numeric_std.ALL;

entity SB_RAM4KNR is

  generic ( 
           TimingChecksOn : boolean := true;
           Xon            : boolean := false;
           MsgOn          : boolean := false;
           
           tipd_RCLKN  : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_RCLKE : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_RE    : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_RADDR : VitalDelayArrayType01(7 downto 0)  := (others => (0 ns, 0 ns));
           tipd_WCLK  : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_WCLKE : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_WE    : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_WADDR : VitalDelayArrayType01(7 downto 0)  := (others => (0 ns, 0 ns));
           tipd_MASK  : VitalDelayArrayType01(15 downto 0)  := (others => (0 ns, 0 ns));
           tipd_WDATA : VitalDelayArrayType01(15 downto 0)  := (others => (0 ns, 0 ns));

           tpd_RCLKN_RDATA : VitalDelayArrayType01(15 downto 0) := (others => (100 ns, 100 ns));

           tsetup_RADDR_RCLKN_negedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           tsetup_RADDR_RCLKN_posedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           tsetup_RCLKE_RCLKN_negedge_posedge : VitalDelayType                   := 0 ns;
           tsetup_RCLKE_RCLKN_posedge_posedge : VitalDelayType                   := 0 ns;
           tsetup_RE_RCLKN_negedge_posedge    : VitalDelayType                   := 0 ns;
           tsetup_RE_RCLKN_posedge_posedge    : VitalDelayType                   := 0 ns;

           tsetup_WADDR_WCLK_negedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           tsetup_WADDR_WCLK_posedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           tsetup_WDATA_WCLK_negedge_posedge : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           tsetup_WDATA_WCLK_posedge_posedge : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           tsetup_WCLKE_WCLK_negedge_posedge : VitalDelayType                   := 0 ns;
           tsetup_WCLKE_WCLK_posedge_posedge : VitalDelayType                   := 0 ns;
           tsetup_WE_WCLK_negedge_posedge    : VitalDelayType                   := 0 ns;
           tsetup_WE_WCLK_posedge_posedge    : VitalDelayType                   := 0 ns;
           tsetup_MASK_WCLK_negedge_posedge  : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           tsetup_MASK_WCLK_posedge_posedge  : VitalDelayArrayType(15 downto 0) := (others => 0 ns);

           thold_RADDR_RCLKN_negedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           thold_RADDR_RCLKN_posedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           thold_RCLKE_RCLKN_negedge_posedge : VitalDelayType                   := 0 ns;
           thold_RCLKE_RCLKN_posedge_posedge : VitalDelayType                   := 0 ns;
           thold_RE_RCLKN_negedge_posedge    : VitalDelayType                   := 0 ns;
           thold_RE_RCLKN_posedge_posedge    : VitalDelayType                   := 0 ns;

           thold_WADDR_WCLK_negedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           thold_WADDR_WCLK_posedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           thold_WDATA_WCLK_negedge_posedge : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           thold_WDATA_WCLK_posedge_posedge : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           thold_WCLKE_WCLK_negedge_posedge : VitalDelayType                   := 0 ns;
           thold_WCLKE_WCLK_posedge_posedge : VitalDelayType                   := 0 ns;
           thold_WE_WCLK_negedge_posedge    : VitalDelayType                   := 0 ns;
           thold_WE_WCLK_posedge_posedge    : VitalDelayType                   := 0 ns;
           thold_MASK_WCLK_negedge_posedge  : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           thold_MASK_WCLK_posedge_posedge  : VitalDelayArrayType(15 downto 0) := (others => 0 ns);

           tpw_RCLKN_negedge : VitalDelayType := 0 ns;
           tpw_RCLKN_posedge : VitalDelayType := 0 ns;
           tpw_WCLK_negedge : VitalDelayType := 0 ns;
           tpw_WCLK_posedge : VitalDelayType := 0 ns;

           trecovery_RCLKN_WCLK_posedge_posedge  : VitalDelayType                   := 0 ns;
           trecovery_RCLKN_WCLK_negedge_posedge  : VitalDelayType                   := 0 ns;
           tremoval_RCLKN_WCLK_posedge_posedge   : VitalDelayType                   := 0 ns;
           tremoval_RCLKN_WCLK_negedge_posedge   : VitalDelayType                   := 0 ns;
           trecovery_WCLK_RCLKN_posedge_posedge  : VitalDelayType                   := 0 ns;
           trecovery_WCLK_RCLKN_negedge_posedge  : VitalDelayType                   := 0 ns;
           tremoval_WCLK_RCLKN_posedge_posedge   : VitalDelayType                   := 0 ns;
           tremoval_WCLK_RCLKN_negedge_posedge   : VitalDelayType                   := 0 ns;


           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 15  downto 0) ;
                RCLKN  : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'L';
                RADDR : in  std_logic_vector( 7  downto 0) ;
                WCLK  : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'L';
                WADDR : in  std_logic_vector( 7  downto 0) ;
                MASK  : in  std_logic_vector( 15  downto 0) ;
                WDATA : in  std_logic_vector( 15  downto 0)
               );
  
  --attribute VITAL_LEVEL0 of SB_RAM4KNR : entity is TRUE;
  
end SB_RAM4KNR;



architecture SB_RAM4KNR_V of SB_RAM4KNR is
    
  --attribute VITAL_LEVEL0 of SB_RAM4KNR_V : architecture is TRUE;

  --signal RDATA_reg : std_logic_vector( 15  downto 0) := (others => '0');

  signal MEM : std_logic_vector(4095 downto 0) ;
  signal Address_Collision_Detected : std_logic ;


  signal RADDR_ipd : std_logic_vector(7 downto 0)  := (others => 'X');
  signal RCLKN_ipd  : std_logic                    := 'X';
  signal RCLKE_ipd : std_logic                    := 'X';
  signal RE_ipd    : std_logic                    := 'X';

  signal WADDR_ipd : std_logic_vector(7 downto 0)  := (others => 'X');
  signal WCLK_ipd  : std_logic                    := 'X';  
  signal WCLKE_ipd : std_logic                    := 'X';
  signal WE_ipd    : std_logic                    := 'X';
  signal MASK_ipd  : std_logic_vector(15 downto 0) := (others => 'X');
  signal WDATA_ipd : std_logic_vector(15 downto 0) := (others => 'X');

  signal RADDR_in : integer range 0 to 255 ;
  signal WADDR_in : integer range 0 to 255 ;

begin

  --RDATA <= RDATA_reg;

---------------------
--  Input Wire Delay
---------------------
  WireDelay : block
  begin
    RADDR_DELAY : for i in 7 downto 0 generate
       VitalWireDelay (RADDR_ipd(i), RADDR(i), tipd_RADDR(i));
    end generate RADDR_DELAY;
    VitalWireDelay (RCLKN_ipd, RCLKN, tipd_RCLKN);
    VitalWireDelay (RCLKE_ipd, RCLKE, tipd_RCLKE);
    VitalWireDelay (RE_ipd, RE, tipd_RE);
    WADDR_DELAY : for i in 7 downto 0 generate
       VitalWireDelay (WADDR_ipd(i), WADDR(i), tipd_WADDR(i));
    end generate WADDR_DELAY;
    VitalWireDelay (WCLK_ipd, WCLK, tipd_WCLK);
    VitalWireDelay (WCLKE_ipd, WCLKE, tipd_WCLKE);
    VitalWireDelay (WE_ipd, WE, tipd_WE);
    MASK_DELAY : for i in 15 downto 0 generate
       VitalWireDelay (MASK_ipd(i), MASK(i), tipd_MASK(i));
    end generate MASK_DELAY;
    WDATA_DELAY : for i in 15 downto 0 generate
       VitalWireDelay (WDATA_ipd(i), WDATA(i), tipd_WDATA(i));
    end generate WDATA_DELAY;
  end block;

  process(RE_ipd,WE_ipd,WADDR_ipd,RADDR_ipd)
      begin
          if ( (WE_ipd = '1')  and (RE_ipd = '1') and ( WADDR_ipd = RADDR_ipd) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;
          assert (not(Address_Collision_Detected = '1'))
            report "Address_Collision"
            severity warning ;         
  end process; 



  VITALReadBehavior : process(RADDR_ipd,RCLKN_ipd,RCLKE_ipd,RE_ipd)
   
       variable Tviol_RADDR0_RCLKN_posedge : std_logic := '0';
       variable Tviol_RADDR1_RCLKN_posedge : std_logic := '0';
       variable Tviol_RADDR2_RCLKN_posedge : std_logic := '0';
       variable Tviol_RADDR3_RCLKN_posedge : std_logic := '0';
       variable Tviol_RADDR4_RCLKN_posedge : std_logic := '0';
       variable Tviol_RADDR5_RCLKN_posedge : std_logic := '0';
       variable Tviol_RADDR6_RCLKN_posedge : std_logic := '0';
       variable Tviol_RADDR7_RCLKN_posedge : std_logic := '0';
       variable Tviol_RCLKE_RCLKN_posedge  : std_logic := '0';
       variable Tviol_RE_RCLKN_posedge     : std_logic := '0';

       variable Tmkr_RADDR0_RCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR1_RCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR2_RCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR3_RCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR4_RCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR5_RCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR6_RCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR7_RCLKN_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RCLKE_RCLKN_posedge  : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RE_RCLKN_posedge     : VitalTimingDataType := VitalTimingDataInit;

       variable PViol_RCLKN : std_logic := '0';

       variable PInfo_RCLKN : VitalPeriodDataType ;

       variable Tviol_WCLK_RCLKN_posedge : std_logic := '0';
       variable Tmkr_WCLK_RCLKN_posedge  : VitalTimingDataType := VitalTimingDataInit ;
       variable Tviol_WCLK_RCLKN_negedge : std_logic := '0';
       variable Tmkr_WCLK_RCLKN_negedge  : VitalTimingDataType := VitalTimingDataInit ;

       variable RDATA_GlitchData0  : VitalGlitchDataType;
       variable RDATA_GlitchData1  : VitalGlitchDataType;
       variable RDATA_GlitchData2  : VitalGlitchDataType;
       variable RDATA_GlitchData3  : VitalGlitchDataType;
       variable RDATA_GlitchData4  : VitalGlitchDataType;
       variable RDATA_GlitchData5  : VitalGlitchDataType;
       variable RDATA_GlitchData6  : VitalGlitchDataType;
       variable RDATA_GlitchData7  : VitalGlitchDataType;
       variable RDATA_GlitchData8  : VitalGlitchDataType;
       variable RDATA_GlitchData9  : VitalGlitchDataType;
       variable RDATA_GlitchData10 : VitalGlitchDataType;
       variable RDATA_GlitchData11 : VitalGlitchDataType;
       variable RDATA_GlitchData12 : VitalGlitchDataType;
       variable RDATA_GlitchData13 : VitalGlitchDataType;
       variable RDATA_GlitchData14 : VitalGlitchDataType;
       variable RDATA_GlitchData15 : VitalGlitchDataType;

       variable Violation     : std_logic  := '0';

       variable temp : std_logic_vector(15 downto 0) := (others => 'X');
       variable RDATA_zd : std_logic_vector(15 downto 0) := (others => 'X');

  begin

  -------------------------
  --  Functionality Section
  -------------------------
    RADDR_in <= conv_integer(RADDR_ipd) ;
  
    if (Violation = '1') then
       RDATA <= (others => 'X') ;
    elsif ( RCLKN_ipd'event and (RCLKN_ipd = '0') and (RCLKE_ipd = '1' or RCLKE_ipd = 'H') and (RE_ipd = '1') ) then
       for i in 0 to 15 loop
         temp(i) := MEM(16*RADDR_in + i ) ;
       end loop ;
    end if ; 

    --RDATA_reg <= temp ;
    RDATA <= temp ;


  ------------------------
  --  Timing Check Section
  ------------------------
    if (TimingChecksOn) then
      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR0_RCLKN_posedge,
        TimingData     => Tmkr_RADDR0_RCLKN_posedge,
        TestSignal     => RADDR_ipd(0),
        TestSignalName => "RADDR(0)",
        TestDelay      => 0 ns,
        RefSignal      => RCLKN_ipd,
        RefSignalName  => "RCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLKN_posedge_posedge(0),
        SetupLow       => tsetup_RADDR_RCLKN_negedge_posedge(0),
        HoldLow        => thold_RADDR_RCLKN_posedge_posedge(0),
        HoldHigh       => thold_RADDR_RCLKN_negedge_posedge(0),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR1_RCLKN_posedge,
        TimingData     => Tmkr_RADDR1_RCLKN_posedge,
        TestSignal     => RADDR_ipd(1),
        TestSignalName => "RADDR(1)",
        TestDelay      => 0 ns,
        RefSignal      => RCLKN_ipd,
        RefSignalName  => "RCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLKN_posedge_posedge(1),
        SetupLow       => tsetup_RADDR_RCLKN_negedge_posedge(1),
        HoldLow        => thold_RADDR_RCLKN_posedge_posedge(1),
        HoldHigh       => thold_RADDR_RCLKN_negedge_posedge(1),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR2_RCLKN_posedge,
        TimingData     => Tmkr_RADDR2_RCLKN_posedge,
        TestSignal     => RADDR_ipd(2),
        TestSignalName => "RADDR(2)",
        TestDelay      => 0 ns,
        RefSignal      => RCLKN_ipd,
        RefSignalName  => "RCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLKN_posedge_posedge(2),
        SetupLow       => tsetup_RADDR_RCLKN_negedge_posedge(2),
        HoldLow        => thold_RADDR_RCLKN_posedge_posedge(2),
        HoldHigh       => thold_RADDR_RCLKN_negedge_posedge(2),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR3_RCLKN_posedge,
        TimingData     => Tmkr_RADDR3_RCLKN_posedge,
        TestSignal     => RADDR_ipd(3),
        TestSignalName => "RADDR(3)",
        TestDelay      => 0 ns,
        RefSignal      => RCLKN_ipd,
        RefSignalName  => "RCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLKN_posedge_posedge(3),
        SetupLow       => tsetup_RADDR_RCLKN_negedge_posedge(3),
        HoldLow        => thold_RADDR_RCLKN_posedge_posedge(3),
        HoldHigh       => thold_RADDR_RCLKN_negedge_posedge(3),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR4_RCLKN_posedge,
        TimingData     => Tmkr_RADDR4_RCLKN_posedge,
        TestSignal     => RADDR_ipd(4),
        TestSignalName => "RADDR(4)",
        TestDelay      => 0 ns,
        RefSignal      => RCLKN_ipd,
        RefSignalName  => "RCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLKN_posedge_posedge(4),
        SetupLow       => tsetup_RADDR_RCLKN_negedge_posedge(4),
        HoldLow        => thold_RADDR_RCLKN_posedge_posedge(4),
        HoldHigh       => thold_RADDR_RCLKN_negedge_posedge(4),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR5_RCLKN_posedge,
        TimingData     => Tmkr_RADDR5_RCLKN_posedge,
        TestSignal     => RADDR_ipd(5),
        TestSignalName => "RADDR(5)",
        TestDelay      => 0 ns,
        RefSignal      => RCLKN_ipd,
        RefSignalName  => "RCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLKN_posedge_posedge(5),
        SetupLow       => tsetup_RADDR_RCLKN_negedge_posedge(5),
        HoldLow        => thold_RADDR_RCLKN_posedge_posedge(5),
        HoldHigh       => thold_RADDR_RCLKN_negedge_posedge(5),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR6_RCLKN_posedge,
        TimingData     => Tmkr_RADDR6_RCLKN_posedge,
        TestSignal     => RADDR_ipd(6),
        TestSignalName => "RADDR(6)",
        TestDelay      => 0 ns,
        RefSignal      => RCLKN_ipd,
        RefSignalName  => "RCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLKN_posedge_posedge(6),
        SetupLow       => tsetup_RADDR_RCLKN_negedge_posedge(6),
        HoldLow        => thold_RADDR_RCLKN_posedge_posedge(6),
        HoldHigh       => thold_RADDR_RCLKN_negedge_posedge(6),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR7_RCLKN_posedge,
        TimingData     => Tmkr_RADDR7_RCLKN_posedge,
        TestSignal     => RADDR_ipd(7),
        TestSignalName => "RADDR(7)",
        TestDelay      => 0 ns,
        RefSignal      => RCLKN_ipd,
        RefSignalName  => "RCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLKN_posedge_posedge(7),
        SetupLow       => tsetup_RADDR_RCLKN_negedge_posedge(7),
        HoldLow        => thold_RADDR_RCLKN_posedge_posedge(7),
        HoldHigh       => thold_RADDR_RCLKN_negedge_posedge(7),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_RCLKE_RCLKN_posedge,
        TimingData     => Tmkr_RCLKE_RCLKN_posedge,
        TestSignal     => RCLKE_ipd,
        TestSignalName => "RCLKE",
        TestDelay      => 0 ns,
        RefSignal      => RCLKN_ipd,
        RefSignalName  => "RCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RCLKE_RCLKN_posedge_posedge,
        SetupLow       => tsetup_RCLKE_RCLKN_negedge_posedge,
        HoldLow        => thold_RCLKE_RCLKN_posedge_posedge,
        HoldHigh       => thold_RCLKE_RCLKN_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_RE_RCLKN_posedge,
        TimingData     => Tmkr_RE_RCLKN_posedge,
        TestSignal     => RCLKN_ipd,
        TestSignalName => "RCLKN",
        TestDelay      => 0 ns,
        RefSignal      => RCLKN_ipd,
        RefSignalName  => "RCLKN",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RE_RCLKN_posedge_posedge,
        SetupLow       => tsetup_RE_RCLKN_negedge_posedge,
        HoldLow        => thold_RE_RCLKN_posedge_posedge,
        HoldHigh       => thold_RE_RCLKN_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
        

      VitalPeriodPulseCheck (
        Violation      => Pviol_RCLKN,
        PeriodData     => PInfo_RCLKN,
        TestSignal     => RCLKN_ipd,
        TestSignalName => "RCLKN",
        TestDelay      => 0 ns,
        Period         => 0 ns,
        PulseWidthHigh => tpw_RCLKN_posedge,
        PulseWidthLow  => tpw_RCLKN_negedge,
        CheckEnabled   => true,
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

     VitalRecoveryRemovalCheck (
       Violation               => Tviol_WCLK_RCLKN_posedge,
       TimingData              => Tmkr_WCLK_RCLKN_posedge,
       TestSignal              => WCLK_ipd,
       TestSignalName          => "WCLK",
       TestDelay               => 0 ns,
       RefSignal               => RCLKN_ipd,
       RefSignalName          => "RCLKN",
       RefDelay                => 0 ns,
       Recovery                => trecovery_WCLK_RCLKN_negedge_posedge,
       Removal                 => tremoval_WCLK_RCLKN_negedge_posedge,
       ActiveLow               => FALSE,
       CheckEnabled            => true,
       RefTransition           => 'R',
       HeaderMsg               => "/SB_RAM4KNR",
       Xon                     => Xon,
       MsgOn                   => MsgOn,
       MsgSeverity             => WARNING);

     VitalRecoveryRemovalCheck (
       Violation               => Tviol_WCLK_RCLKN_negedge,
       TimingData              => Tmkr_WCLK_RCLKN_negedge,
       TestSignal              => WCLK_ipd,
       TestSignalName          => "WCLK",
       TestDelay               => 0 ns,
       RefSignal               => RCLKN_ipd,
       RefSignalName          => "RCLKN",
       RefDelay                => 0 ns,
       Recovery                => trecovery_WCLK_RCLKN_posedge_posedge,
       Removal                 => tremoval_WCLK_RCLKN_posedge_posedge,
       ActiveLow               => FALSE,
       CheckEnabled            => true,
       RefTransition           => 'R',
       HeaderMsg               => "/SB_RAM4KNR",
       Xon                     => Xon,
       MsgOn                   => MsgOn,
       MsgSeverity             => WARNING);


    end if ;

    Violation  := Pviol_RCLKN or
                  Tviol_RADDR0_RCLKN_posedge or
                  Tviol_RADDR1_RCLKN_posedge or
                  Tviol_RADDR2_RCLKN_posedge or
                  Tviol_RADDR3_RCLKN_posedge or
                  Tviol_RADDR4_RCLKN_posedge or
                  Tviol_RADDR5_RCLKN_posedge or
                  Tviol_RADDR6_RCLKN_posedge or
                  Tviol_RADDR7_RCLKN_posedge or
                  Tviol_RCLKE_RCLKN_posedge or
                  Tviol_RE_RCLKN_posedge or
                  Tviol_WCLK_RCLKN_posedge or
                  Tviol_WCLK_RCLKN_negedge;

    RDATA_zd(0) := Violation xor RDATA_zd(0) ;
    RDATA_zd(1) := Violation xor RDATA_zd(1) ;
    RDATA_zd(2) := Violation xor RDATA_zd(2) ;
    RDATA_zd(3) := Violation xor RDATA_zd(3) ;
    RDATA_zd(4) := Violation xor RDATA_zd(4) ;
    RDATA_zd(5) := Violation xor RDATA_zd(5) ;
    RDATA_zd(6) := Violation xor RDATA_zd(6) ;
    RDATA_zd(7) := Violation xor RDATA_zd(7) ;
    RDATA_zd(8) := Violation xor RDATA_zd(8) ;
    RDATA_zd(9) := Violation xor RDATA_zd(9) ;
    RDATA_zd(10) := Violation xor RDATA_zd(10) ;
    RDATA_zd(11) := Violation xor RDATA_zd(11) ;
    RDATA_zd(12) := Violation xor RDATA_zd(12) ;
    RDATA_zd(13) := Violation xor RDATA_zd(13) ;
    RDATA_zd(14) := Violation xor RDATA_zd(14) ;
    RDATA_zd(15) := Violation xor RDATA_zd(15) ;
    
    
    
    
    
  ----------------------
  --  Path Delay Section
  ----------------------
    VitalPathDelay01 (
      OutSignal     => RDATA(0),
      GlitchData    => RDATA_GlitchData0,
      OutSignalName => "RDATA(0)",
      OutTemp       => RDATA_zd(0),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(0), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(1),
      GlitchData    => RDATA_GlitchData1,
      OutSignalName => "RDATA(1)",
      OutTemp       => RDATA_zd(1),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(1), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(2),
      GlitchData    => RDATA_GlitchData2,
      OutSignalName => "RDATA(2)",
      OutTemp       => RDATA_zd(2),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(2), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(3),
      GlitchData    => RDATA_GlitchData3,
      OutSignalName => "RDATA(3)",
      OutTemp       => RDATA_zd(3),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(3), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(4),
      GlitchData    => RDATA_GlitchData4,
      OutSignalName => "RDATA(4)",
      OutTemp       => RDATA_zd(4),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(4), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(5),
      GlitchData    => RDATA_GlitchData5,
      OutSignalName => "RDATA(5)",
      OutTemp       => RDATA_zd(5),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(5), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(6),
      GlitchData    => RDATA_GlitchData6,
      OutSignalName => "RDATA(6)",
      OutTemp       => RDATA_zd(6),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(6), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(7),
      GlitchData    => RDATA_GlitchData7,
      OutSignalName => "RDATA(7)",
      OutTemp       => RDATA_zd(7),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(7), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(8),
      GlitchData    => RDATA_GlitchData8,
      OutSignalName => "RDATA(8)",
      OutTemp       => RDATA_zd(8),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(8), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(9),
      GlitchData    => RDATA_GlitchData9,
      OutSignalName => "RDATA(9)",
      OutTemp       => RDATA_zd(9),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(9), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(10),
      GlitchData    => RDATA_GlitchData10,
      OutSignalName => "RDATA(10)",
      OutTemp       => RDATA_zd(10),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(10), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(11),
      GlitchData    => RDATA_GlitchData11,
      OutSignalName => "RDATA(11)",
      OutTemp       => RDATA_zd(11),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(11), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(12),
      GlitchData    => RDATA_GlitchData12,
      OutSignalName => "RDATA(12)",
      OutTemp       => RDATA_zd(12),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(12), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(13),
      GlitchData    => RDATA_GlitchData13,
      OutSignalName => "RDATA(13)",
      OutTemp       => RDATA_zd(13),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(13), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(14),
      GlitchData    => RDATA_GlitchData14,
      OutSignalName => "RDATA(14)",
      OutTemp       => RDATA_zd(14),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(14), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(15),
      GlitchData    => RDATA_GlitchData15,
      OutSignalName => "RDATA(15)",
      OutTemp       => RDATA_zd(15),
      Paths         => (0 => (RCLKN_ipd'last_event, tpd_RCLKN_RDATA(15), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);




  end process VITALReadBehavior;

  VITALWriteBehavior : process(WADDR_ipd,WCLK_ipd,WCLKE_ipd,WE_ipd)

       variable Tviol_WADDR0_WCLK_posedge : std_logic := '0';
       variable Tviol_WADDR1_WCLK_posedge : std_logic := '0';
       variable Tviol_WADDR2_WCLK_posedge : std_logic := '0';
       variable Tviol_WADDR3_WCLK_posedge : std_logic := '0';
       variable Tviol_WADDR4_WCLK_posedge : std_logic := '0';
       variable Tviol_WADDR5_WCLK_posedge : std_logic := '0';
       variable Tviol_WADDR6_WCLK_posedge : std_logic := '0';
       variable Tviol_WADDR7_WCLK_posedge : std_logic := '0';
       variable Tviol_WCLKE_WCLK_posedge  : std_logic := '0';
       variable Tviol_WE_WCLK_posedge     : std_logic := '0';
       variable Tviol_WDATA0_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA1_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA2_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA3_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA4_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA5_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA6_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA7_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA8_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA9_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA10_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA11_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA12_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA13_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA14_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA15_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK0_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK1_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK2_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK3_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK4_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK5_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK6_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK7_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK8_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK9_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK10_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK11_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK12_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK13_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK14_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK15_WCLK_posedge : std_logic := '0';


       variable Tmkr_WADDR0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR5_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR6_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR7_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WCLKE_WCLK_posedge  : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WE_WCLK_posedge     : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA5_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA6_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA7_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA8_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA9_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA10_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA11_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA12_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA13_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA14_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA15_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK5_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK6_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK7_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK8_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK9_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK10_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK11_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK12_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK13_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK14_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK15_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;

       variable PViol_WCLK : std_logic := '0';

       variable PInfo_WCLK : VitalPeriodDataType := VitalPeriodDataInit;

       variable Tviol_RCLKN_WCLK_posedge : std_logic := '0';
       variable Tmkr_RCLKN_WCLK_posedge  : VitalTimingDataType := VitalTimingDataInit;
       variable Tviol_RCLKN_WCLK_negedge : std_logic := '0';
       variable Tmkr_RCLKN_WCLK_negedge  : VitalTimingDataType := VitalTimingDataInit;


       variable Violation     : std_logic  := '0';

       variable MEM_temp : std_logic_vector(4095 downto 0) := To_StdLogicVector(INIT_F) &
                                                              To_StdLogicVector(INIT_E) &
                                                              To_StdLogicVector(INIT_D) &
                                                              To_StdLogicVector(INIT_C) &
                                                              To_StdLogicVector(INIT_B) &
                                                              To_StdLogicVector(INIT_A) &
                                                              To_StdLogicVector(INIT_9) &
                                                              To_StdLogicVector(INIT_8) &
                                                              To_StdLogicVector(INIT_7) &
                                                              To_StdLogicVector(INIT_6) &
                                                              To_StdLogicVector(INIT_5) &
                                                              To_StdLogicVector(INIT_4) &
                                                              To_StdLogicVector(INIT_3) &
                                                              To_StdLogicVector(INIT_2) &
                                                              To_StdLogicVector(INIT_1) &
                                                              To_StdLogicVector(INIT_0);
       
  begin

    Violation  := Pviol_WCLK or
                  Tviol_WADDR0_WCLK_posedge or
                  Tviol_WADDR1_WCLK_posedge or
                  Tviol_WADDR2_WCLK_posedge or
                  Tviol_WADDR3_WCLK_posedge or
                  Tviol_WADDR4_WCLK_posedge or
                  Tviol_WADDR5_WCLK_posedge or
                  Tviol_WADDR6_WCLK_posedge or
                  Tviol_WADDR7_WCLK_posedge or
                  Tviol_WCLKE_WCLK_posedge or
                  Tviol_WE_WCLK_posedge or
                  Tviol_WDATA0_WCLK_posedge or
                  Tviol_WDATA1_WCLK_posedge or
                  Tviol_WDATA2_WCLK_posedge or
                  Tviol_WDATA3_WCLK_posedge or
                  Tviol_WDATA4_WCLK_posedge or
                  Tviol_WDATA5_WCLK_posedge or
                  Tviol_WDATA6_WCLK_posedge or
                  Tviol_WDATA7_WCLK_posedge or
                  Tviol_WDATA8_WCLK_posedge or
                  Tviol_WDATA9_WCLK_posedge or
                  Tviol_WDATA10_WCLK_posedge or
                  Tviol_WDATA11_WCLK_posedge or
                  Tviol_WDATA12_WCLK_posedge or
                  Tviol_WDATA13_WCLK_posedge or
                  Tviol_WDATA14_WCLK_posedge or
                  Tviol_WDATA15_WCLK_posedge or
                  Tviol_MASK0_WCLK_posedge or
                  Tviol_MASK1_WCLK_posedge or
                  Tviol_MASK2_WCLK_posedge or
                  Tviol_MASK3_WCLK_posedge or
                  Tviol_MASK4_WCLK_posedge or
                  Tviol_MASK5_WCLK_posedge or
                  Tviol_MASK6_WCLK_posedge or
                  Tviol_MASK7_WCLK_posedge or
                  Tviol_MASK8_WCLK_posedge or
                  Tviol_MASK9_WCLK_posedge or
                  Tviol_MASK10_WCLK_posedge or
                  Tviol_MASK11_WCLK_posedge or
                  Tviol_MASK12_WCLK_posedge or
                  Tviol_MASK13_WCLK_posedge or
                  Tviol_MASK14_WCLK_posedge or
                  Tviol_MASK15_WCLK_posedge or
                  Tviol_RCLKN_WCLK_posedge or
                  Tviol_RCLKN_WCLK_negedge;
 
-------------------------
--  Functionality Section
-------------------------

    WADDR_in <= conv_integer(WADDR_ipd) ;
  
    if (Violation = '1') then
       MEM <= (others => 'X') ;
    elsif ( WCLK_ipd'event and (WCLK_ipd = '1') and (WCLKE_ipd = '1' or WCLKE_ipd = 'H') and (WE_ipd = '1') ) then
       for i in 0 to 15 loop
         if (MASK(i) = '0') then
            MEM_temp(16*WADDR_in + i ) := WDATA_ipd(i) ;
         end if ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;

------------------------
--  Timing Check Section
------------------------
    if (TimingChecksOn) then
      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR0_WCLK_posedge,
        TimingData     => Tmkr_WADDR0_WCLK_posedge,
        TestSignal     => WADDR_ipd(0),
        TestSignalName => "WADDR(0)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(0),
        SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(0),
        HoldLow        => thold_WADDR_WCLK_posedge_posedge(0),
        HoldHigh       => thold_WADDR_WCLK_negedge_posedge(0),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR1_WCLK_posedge,
        TimingData     => Tmkr_WADDR1_WCLK_posedge,
        TestSignal     => WADDR_ipd(1),
        TestSignalName => "WADDR(1)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(1),
        SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(1),
        HoldLow        => thold_WADDR_WCLK_posedge_posedge(1),
        HoldHigh       => thold_WADDR_WCLK_negedge_posedge(1),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR2_WCLK_posedge,
        TimingData     => Tmkr_WADDR2_WCLK_posedge,
        TestSignal     => WADDR_ipd(2),
        TestSignalName => "WADDR(2)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(2),
        SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(2),
        HoldLow        => thold_WADDR_WCLK_posedge_posedge(2),
        HoldHigh       => thold_WADDR_WCLK_negedge_posedge(2),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR3_WCLK_posedge,
        TimingData     => Tmkr_WADDR3_WCLK_posedge,
        TestSignal     => WADDR_ipd(3),
        TestSignalName => "WADDR(3)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(3),
        SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(3),
        HoldLow        => thold_WADDR_WCLK_posedge_posedge(3),
        HoldHigh       => thold_WADDR_WCLK_negedge_posedge(3),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR4_WCLK_posedge,
        TimingData     => Tmkr_WADDR4_WCLK_posedge,
        TestSignal     => WADDR_ipd(4),
        TestSignalName => "WADDR(4)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(4),
        SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(4),
        HoldLow        => thold_WADDR_WCLK_posedge_posedge(4),
        HoldHigh       => thold_WADDR_WCLK_negedge_posedge(4),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR5_WCLK_posedge,
        TimingData     => Tmkr_WADDR5_WCLK_posedge,
        TestSignal     => WADDR_ipd(5),
        TestSignalName => "WADDR(5)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(5),
        SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(5),
        HoldLow        => thold_WADDR_WCLK_posedge_posedge(5),
        HoldHigh       => thold_WADDR_WCLK_negedge_posedge(5),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR6_WCLK_posedge,
        TimingData     => Tmkr_WADDR6_WCLK_posedge,
        TestSignal     => WADDR_ipd(6),
        TestSignalName => "WADDR(6)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(6),
        SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(6),
        HoldLow        => thold_WADDR_WCLK_posedge_posedge(6),
        HoldHigh       => thold_WADDR_WCLK_negedge_posedge(6),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR7_WCLK_posedge,
        TimingData     => Tmkr_WADDR7_WCLK_posedge,
        TestSignal     => WADDR_ipd(7),
        TestSignalName => "WADDR(7)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(7),
        SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(7),
        HoldLow        => thold_WADDR_WCLK_posedge_posedge(7),
        HoldHigh       => thold_WADDR_WCLK_negedge_posedge(7),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WCLKE_WCLK_posedge,
        TimingData     => Tmkr_WCLKE_WCLK_posedge,
        TestSignal     => WCLKE_ipd,
        TestSignalName => "WCLKE",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WCLKE_WCLK_posedge_posedge,
        SetupLow       => tsetup_WCLKE_WCLK_negedge_posedge,
        HoldLow        => thold_WCLKE_WCLK_posedge_posedge,
        HoldHigh       => thold_WCLKE_WCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WE_WCLK_posedge,
        TimingData     => Tmkr_WE_WCLK_posedge,
        TestSignal     => WCLK_ipd,
        TestSignalName => "WCLK",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WE_WCLK_posedge_posedge,
        SetupLow       => tsetup_WE_WCLK_negedge_posedge,
        HoldLow        => thold_WE_WCLK_posedge_posedge,
        HoldHigh       => thold_WE_WCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
       VitalSetupHoldCheck (
        Violation      => Tviol_WDATA0_WCLK_posedge,
        TimingData     => Tmkr_WDATA0_WCLK_posedge,
        TestSignal     => WDATA_ipd(0),
        TestSignalName => "WDATA(0)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(0),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(0),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(0),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(0),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA1_WCLK_posedge,
        TimingData     => Tmkr_WDATA1_WCLK_posedge,
        TestSignal     => WDATA_ipd(1),
        TestSignalName => "WDATA(1)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(1),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(1),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(1),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(1),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA2_WCLK_posedge,
        TimingData     => Tmkr_WDATA2_WCLK_posedge,
        TestSignal     => WDATA_ipd(2),
        TestSignalName => "WDATA(2)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(2),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(2),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(2),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(2),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA3_WCLK_posedge,
        TimingData     => Tmkr_WDATA3_WCLK_posedge,
        TestSignal     => WDATA_ipd(3),
        TestSignalName => "WDATA(3)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(3),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(3),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(3),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(3),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA4_WCLK_posedge,
        TimingData     => Tmkr_WDATA4_WCLK_posedge,
        TestSignal     => WDATA_ipd(4),
        TestSignalName => "WDATA(4)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(4),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(4),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(4),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(4),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA5_WCLK_posedge,
        TimingData     => Tmkr_WDATA5_WCLK_posedge,
        TestSignal     => WDATA_ipd(5),
        TestSignalName => "WDATA(5)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(5),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(5),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(5),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(5),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA6_WCLK_posedge,
        TimingData     => Tmkr_WDATA6_WCLK_posedge,
        TestSignal     => WDATA_ipd(6),
        TestSignalName => "WDATA(6)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(6),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(6),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(6),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(6),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA7_WCLK_posedge,
        TimingData     => Tmkr_WDATA7_WCLK_posedge,
        TestSignal     => WDATA_ipd(7),
        TestSignalName => "WDATA(7)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(7),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(7),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(7),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(7),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

       VitalSetupHoldCheck (
        Violation      => Tviol_WDATA8_WCLK_posedge,
        TimingData     => Tmkr_WDATA8_WCLK_posedge,
        TestSignal     => WDATA_ipd(8),
        TestSignalName => "WDATA(8)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(8),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(8),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(8),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(8),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA9_WCLK_posedge,
        TimingData     => Tmkr_WDATA9_WCLK_posedge,
        TestSignal     => WDATA_ipd(9),
        TestSignalName => "WDATA(9)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(9),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(9),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(9),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(9),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA10_WCLK_posedge,
        TimingData     => Tmkr_WDATA10_WCLK_posedge,
        TestSignal     => WDATA_ipd(10),
        TestSignalName => "WDATA(10)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(10),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(10),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(10),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(10),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA11_WCLK_posedge,
        TimingData     => Tmkr_WDATA11_WCLK_posedge,
        TestSignal     => WDATA_ipd(11),
        TestSignalName => "WDATA(11)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(11),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(11),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(11),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(11),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA12_WCLK_posedge,
        TimingData     => Tmkr_WDATA12_WCLK_posedge,
        TestSignal     => WDATA_ipd(12),
        TestSignalName => "WDATA(12)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(12),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(12),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(12),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(12),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA13_WCLK_posedge,
        TimingData     => Tmkr_WDATA13_WCLK_posedge,
        TestSignal     => WDATA_ipd(13),
        TestSignalName => "WDATA(13)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(13),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(13),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(13),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(13),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA14_WCLK_posedge,
        TimingData     => Tmkr_WDATA14_WCLK_posedge,
        TestSignal     => WDATA_ipd(14),
        TestSignalName => "WDATA(14)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(14),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(14),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(14),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(14),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA15_WCLK_posedge,
        TimingData     => Tmkr_WDATA15_WCLK_posedge,
        TestSignal     => WDATA_ipd(15),
        TestSignalName => "WDATA(15)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(15),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(15),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(15),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(15),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

       VitalSetupHoldCheck (
        Violation      => Tviol_MASK0_WCLK_posedge,
        TimingData     => Tmkr_MASK0_WCLK_posedge,
        TestSignal     => MASK_ipd(0),
        TestSignalName => "MASK(0)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(0),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(0),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(0),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(0),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK1_WCLK_posedge,
        TimingData     => Tmkr_MASK1_WCLK_posedge,
        TestSignal     => MASK_ipd(1),
        TestSignalName => "MASK(1)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(1),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(1),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(1),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(1),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK2_WCLK_posedge,
        TimingData     => Tmkr_MASK2_WCLK_posedge,
        TestSignal     => MASK_ipd(2),
        TestSignalName => "MASK(2)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(2),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(2),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(2),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(2),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK3_WCLK_posedge,
        TimingData     => Tmkr_MASK3_WCLK_posedge,
        TestSignal     => MASK_ipd(3),
        TestSignalName => "MASK(3)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(3),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(3),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(3),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(3),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK4_WCLK_posedge,
        TimingData     => Tmkr_MASK4_WCLK_posedge,
        TestSignal     => MASK_ipd(4),
        TestSignalName => "MASK(4)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(4),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(4),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(4),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(4),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_MASK5_WCLK_posedge,
        TimingData     => Tmkr_MASK5_WCLK_posedge,
        TestSignal     => MASK_ipd(5),
        TestSignalName => "MASK(5)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(5),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(5),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(5),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(5),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_MASK6_WCLK_posedge,
        TimingData     => Tmkr_MASK6_WCLK_posedge,
        TestSignal     => MASK_ipd(6),
        TestSignalName => "MASK(6)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(6),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(6),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(6),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(6),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_MASK7_WCLK_posedge,
        TimingData     => Tmkr_MASK7_WCLK_posedge,
        TestSignal     => MASK_ipd(7),
        TestSignalName => "MASK(7)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(7),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(7),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(7),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(7),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

       VitalSetupHoldCheck (
        Violation      => Tviol_MASK8_WCLK_posedge,
        TimingData     => Tmkr_MASK8_WCLK_posedge,
        TestSignal     => MASK_ipd(8),
        TestSignalName => "MASK(8)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(8),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(8),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(8),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(8),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK9_WCLK_posedge,
        TimingData     => Tmkr_MASK9_WCLK_posedge,
        TestSignal     => MASK_ipd(9),
        TestSignalName => "MASK(9)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(9),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(9),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(9),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(9),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK10_WCLK_posedge,
        TimingData     => Tmkr_MASK10_WCLK_posedge,
        TestSignal     => MASK_ipd(10),
        TestSignalName => "MASK(10)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(10),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(10),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(10),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(10),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK11_WCLK_posedge,
        TimingData     => Tmkr_MASK11_WCLK_posedge,
        TestSignal     => MASK_ipd(11),
        TestSignalName => "MASK(11)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(11),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(11),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(11),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(11),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK12_WCLK_posedge,
        TimingData     => Tmkr_MASK12_WCLK_posedge,
        TestSignal     => MASK_ipd(12),
        TestSignalName => "MASK(12)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(12),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(12),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(12),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(12),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_MASK13_WCLK_posedge,
        TimingData     => Tmkr_MASK13_WCLK_posedge,
        TestSignal     => MASK_ipd(13),
        TestSignalName => "MASK(13)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(13),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(13),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(13),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(13),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_MASK14_WCLK_posedge,
        TimingData     => Tmkr_MASK14_WCLK_posedge,
        TestSignal     => MASK_ipd(14),
        TestSignalName => "MASK(14)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(14),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(14),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(14),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(14),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_MASK15_WCLK_posedge,
        TimingData     => Tmkr_MASK15_WCLK_posedge,
        TestSignal     => MASK_ipd(15),
        TestSignalName => "MASK(15)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(15),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(15),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(15),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(15),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
   

      VitalPeriodPulseCheck (
        Violation      => Pviol_WCLK,
        PeriodData     => PInfo_WCLK,
        TestSignal     => WCLK_ipd,
        TestSignalName => "WCLK",
        TestDelay      => 0 ns,
        Period         => 0 ns,
        PulseWidthHigh => tpw_WCLK_posedge,
        PulseWidthLow  => tpw_WCLK_negedge,
        CheckEnabled   => true,
        HeaderMsg      => "/SB_RAM4KNR",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);


     VitalRecoveryRemovalCheck (
       Violation               => Tviol_RCLKN_WCLK_posedge,
       TimingData              => Tmkr_RCLKN_WCLK_posedge,
       TestSignal              => RCLKN_ipd,
       TestSignalName          => "RCLKN",
       TestDelay               => 0 ns,
       RefSignal               => WCLK_ipd,
       RefSignalName          => "WCLK",
       RefDelay                => 0 ns,
       Recovery                => trecovery_RCLKN_WCLK_negedge_posedge,
       Removal                 => tremoval_RCLKN_WCLK_negedge_posedge,
       ActiveLow               => FALSE,
       CheckEnabled            => true,
       RefTransition           => 'R',
       HeaderMsg               => "/SB_RAM4KNR",
       Xon                     => Xon,
       MsgOn                   => MsgOn,
       MsgSeverity             => WARNING);

     VitalRecoveryRemovalCheck (
       Violation               => Tviol_RCLKN_WCLK_negedge,
       TimingData              => Tmkr_RCLKN_WCLK_negedge,
       TestSignal              => RCLKN_ipd,
       TestSignalName          => "RCLKN",
       TestDelay               => 0 ns,
       RefSignal               => WCLK_ipd,
       RefSignalName          => "WCLK",
       RefDelay                => 0 ns,
       Recovery                => trecovery_RCLKN_WCLK_posedge_posedge,
       Removal                 => tremoval_WCLK_RCLKN_posedge_posedge,
       ActiveLow               => FALSE,
       CheckEnabled            => true,
       RefTransition           => 'R',
       HeaderMsg               => "/SB_RAM4KNR",
       Xon                     => Xon,
       MsgOn                   => MsgOn,
       MsgSeverity             => WARNING);


    end if ;


  end process VITALWriteBehavior;


end SB_RAM4KNR_V;



----- CELL SB_RAM4K -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
use IEEE.VITAL_Timing.all; 
USE IEEE.numeric_std.ALL;

entity SB_RAM4K is

  generic ( 
           TimingChecksOn : boolean := true;
           Xon            : boolean := false;
           MsgOn          : boolean := false;
           
           tipd_RCLK  : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_RCLKE : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_RE    : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_RADDR : VitalDelayArrayType01(7 downto 0)  := (others => (0 ns, 0 ns));
           tipd_WCLK  : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_WCLKE : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_WE    : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_WADDR : VitalDelayArrayType01(7 downto 0)  := (others => (0 ns, 0 ns));
           tipd_MASK  : VitalDelayArrayType01(15 downto 0)  := (others => (0 ns, 0 ns));
           tipd_WDATA : VitalDelayArrayType01(15 downto 0)  := (others => (0 ns, 0 ns));

           tpd_RCLK_RDATA : VitalDelayArrayType01(15 downto 0) := (others => (100 ns, 100 ns));
           tpd_RCLK_RDATA_posedge : VitalDelayArrayType01(15 downto 0) := (others => (100 ns, 100 ns));

           tsetup_RADDR_RCLK_negedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           tsetup_RADDR_RCLK_posedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           tsetup_RCLKE_RCLK_negedge_posedge : VitalDelayType                   := 0 ns;
           tsetup_RCLKE_RCLK_posedge_posedge : VitalDelayType                   := 0 ns;
           tsetup_RE_RCLK_negedge_posedge    : VitalDelayType                   := 0 ns;
           tsetup_RE_RCLK_posedge_posedge    : VitalDelayType                   := 0 ns;

           tsetup_WADDR_WCLK_negedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           tsetup_WADDR_WCLK_posedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           tsetup_WDATA_WCLK_negedge_posedge : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           tsetup_WDATA_WCLK_posedge_posedge : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           tsetup_WCLKE_WCLK_negedge_posedge : VitalDelayType                   := 0 ns;
           tsetup_WCLKE_WCLK_posedge_posedge : VitalDelayType                   := 0 ns;
           tsetup_WE_WCLK_negedge_posedge    : VitalDelayType                   := 0 ns;
           tsetup_WE_WCLK_posedge_posedge    : VitalDelayType                   := 0 ns;
           tsetup_MASK_WCLK_negedge_posedge  : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           tsetup_MASK_WCLK_posedge_posedge  : VitalDelayArrayType(15 downto 0) := (others => 0 ns);

           thold_RADDR_RCLK_negedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           thold_RADDR_RCLK_posedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           thold_RCLKE_RCLK_negedge_posedge : VitalDelayType                   := 0 ns;
           thold_RCLKE_RCLK_posedge_posedge : VitalDelayType                   := 0 ns;
           thold_RE_RCLK_negedge_posedge    : VitalDelayType                   := 0 ns;
           thold_RE_RCLK_posedge_posedge    : VitalDelayType                   := 0 ns;

           thold_WADDR_WCLK_negedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           thold_WADDR_WCLK_posedge_posedge : VitalDelayArrayType(7 downto 0)  := (others => 0 ns);
           thold_WDATA_WCLK_negedge_posedge : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           thold_WDATA_WCLK_posedge_posedge : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           thold_WCLKE_WCLK_negedge_posedge : VitalDelayType                   := 0 ns;
           thold_WCLKE_WCLK_posedge_posedge : VitalDelayType                   := 0 ns;
           thold_WE_WCLK_negedge_posedge    : VitalDelayType                   := 0 ns;
           thold_WE_WCLK_posedge_posedge    : VitalDelayType                   := 0 ns;
           thold_MASK_WCLK_negedge_posedge  : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           thold_MASK_WCLK_posedge_posedge  : VitalDelayArrayType(15 downto 0) := (others => 0 ns);

           tpw_RCLK_negedge : VitalDelayType := 0 ns;
           tpw_RCLK_posedge : VitalDelayType := 0 ns;
           tpw_WCLK_negedge : VitalDelayType := 0 ns;
           tpw_WCLK_posedge : VitalDelayType := 0 ns;


           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 15  downto 0) ;
                RCLK  : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'L';
                RADDR : in  std_logic_vector( 7  downto 0) ;
                WCLK  : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'L';
                WADDR : in  std_logic_vector( 7  downto 0) ;
                MASK  : in  std_logic_vector( 15  downto 0) ;
                WDATA : in  std_logic_vector( 15  downto 0)
               );
  
  --attribute VITAL_LEVEL0 of SB_RAM4K : entity is TRUE;
  
end SB_RAM4K;



architecture SB_RAM4K_V of SB_RAM4K is
    
  --attribute VITAL_LEVEL0 of SB_RAM4K_V : architecture is TRUE;

  --signal RDATA_reg : std_logic_vector( 15  downto 0) := (others => '0');


  signal MEM : std_logic_vector(4095 downto 0) ;
  signal Address_Collision_Detected : std_logic ;


  signal RADDR_ipd : std_logic_vector(7 downto 0)  := (others => 'X');   
  signal RCLK_ipd  : std_logic                    := 'X';
  signal RCLKE_ipd : std_logic                    := 'X';
  signal RE_ipd    : std_logic                    := 'X';

  signal WADDR_ipd : std_logic_vector(7 downto 0)  := (others => 'X');
  signal WCLK_ipd  : std_logic                    := 'X';  
  signal WCLKE_ipd : std_logic                    := 'X';
  signal WE_ipd    : std_logic                    := 'X';
  signal MASK_ipd  : std_logic_vector(15 downto 0) := (others => 'X');
  signal WDATA_ipd : std_logic_vector(15 downto 0) := (others => 'X');

  signal RADDR_in : integer range 0 to 255 ;
  signal WADDR_in : integer range 0 to 255 ;

begin

  --RDATA <= RDATA_reg;

---------------------
--  Input Wire Delay
---------------------
  WireDelay : block
  begin
    RADDR_DELAY : for i in 7 downto 0 generate
       VitalWireDelay (RADDR_ipd(i), RADDR(i), tipd_RADDR(i));
    end generate RADDR_DELAY;
    VitalWireDelay (RCLK_ipd, RCLK, tipd_RCLK);
    VitalWireDelay (RCLKE_ipd, RCLKE, tipd_RCLKE);
    VitalWireDelay (RE_ipd, RE, tipd_RE);
    WADDR_DELAY : for i in 7 downto 0 generate
       VitalWireDelay (WADDR_ipd(i), WADDR(i), tipd_WADDR(i));
    end generate WADDR_DELAY;
    VitalWireDelay (WCLK_ipd, WCLK, tipd_WCLK);
    VitalWireDelay (WCLKE_ipd, WCLKE, tipd_WCLKE);
    VitalWireDelay (WE_ipd, WE, tipd_WE);
    MASK_DELAY : for i in 15 downto 0 generate
       VitalWireDelay (MASK_ipd(i), MASK(i), tipd_MASK(i));
    end generate MASK_DELAY;
    WDATA_DELAY : for i in 15 downto 0 generate
       VitalWireDelay (WDATA_ipd(i), WDATA(i), tipd_WDATA(i));
    end generate WDATA_DELAY;
  end block;

  process(RE_ipd,WE_ipd,WADDR_ipd,RADDR_ipd)
      begin
          if ( (WE_ipd = '1')  and (RE_ipd = '1') and ( WADDR_ipd = RADDR_ipd) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;
          assert (not(Address_Collision_Detected = '1'))
            report "Address_Collision"
            severity warning ;         
  end process; 



  VITALReadBehavior : process(RADDR_ipd,RCLK_ipd,RCLKE_ipd,RE_ipd)
   
       variable Tviol_RADDR0_RCLK_posedge : std_logic := '0';
       variable Tviol_RADDR1_RCLK_posedge : std_logic := '0';
       variable Tviol_RADDR2_RCLK_posedge : std_logic := '0';
       variable Tviol_RADDR3_RCLK_posedge : std_logic := '0';
       variable Tviol_RADDR4_RCLK_posedge : std_logic := '0';
       variable Tviol_RADDR5_RCLK_posedge : std_logic := '0';
       variable Tviol_RADDR6_RCLK_posedge : std_logic := '0';
       variable Tviol_RADDR7_RCLK_posedge : std_logic := '0';
       variable Tviol_RCLKE_RCLK_posedge  : std_logic := '0';
       variable Tviol_RE_RCLK_posedge     : std_logic := '0';

       variable Tmkr_RADDR0_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR1_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR2_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR3_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR4_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR5_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR6_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR7_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RCLKE_RCLK_posedge  : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RE_RCLK_posedge     : VitalTimingDataType := VitalTimingDataInit;

       variable PViol_RCLK : std_logic := '0';

       variable PInfo_RCLK : VitalPeriodDataType ;

       variable RDATA_GlitchData0  : VitalGlitchDataType;
       variable RDATA_GlitchData1  : VitalGlitchDataType;
       variable RDATA_GlitchData2  : VitalGlitchDataType;
       variable RDATA_GlitchData3  : VitalGlitchDataType;
       variable RDATA_GlitchData4  : VitalGlitchDataType;
       variable RDATA_GlitchData5  : VitalGlitchDataType;
       variable RDATA_GlitchData6  : VitalGlitchDataType;
       variable RDATA_GlitchData7  : VitalGlitchDataType;
       variable RDATA_GlitchData8  : VitalGlitchDataType;
       variable RDATA_GlitchData9  : VitalGlitchDataType;
       variable RDATA_GlitchData10 : VitalGlitchDataType;
       variable RDATA_GlitchData11 : VitalGlitchDataType;
       variable RDATA_GlitchData12 : VitalGlitchDataType;
       variable RDATA_GlitchData13 : VitalGlitchDataType;
       variable RDATA_GlitchData14 : VitalGlitchDataType;
       variable RDATA_GlitchData15 : VitalGlitchDataType;

       variable Violation     : std_logic  := '0';

       variable temp : std_logic_vector(15 downto 0) := (others => 'X');   --X 
       variable RDATA_zd : std_logic_vector(15 downto 0) := (others => 'X'); --X 

  begin

  -------------------------
  --  Functionality Section
  -------------------------
    RADDR_in <= conv_integer(RADDR_ipd) ;
  
    if (Violation = '1') then
       RDATA <= (others => 'X') ;
    elsif ( RCLK_ipd'event and (RCLK_ipd = '1') and (RCLKE_ipd = '1' or RCLKE_ipd = 'H') and (RE_ipd = '1') ) then
       for i in 0 to 15 loop
         temp(i) := MEM(16*RADDR_in + i ) ;
       end loop ;
    end if ; 

    --RDATA_reg <= temp ;
    RDATA <= temp;


  ------------------------
  --  Timing Check Section
  ------------------------
    if (TimingChecksOn) then
      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR0_RCLK_posedge,
        TimingData     => Tmkr_RADDR0_RCLK_posedge,
        TestSignal     => RADDR_ipd(0),
        TestSignalName => "RADDR(0)",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(0),
        SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(0),
        HoldLow        => thold_RADDR_RCLK_posedge_posedge(0),
        HoldHigh       => thold_RADDR_RCLK_negedge_posedge(0),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR1_RCLK_posedge,
        TimingData     => Tmkr_RADDR1_RCLK_posedge,
        TestSignal     => RADDR_ipd(1),
        TestSignalName => "RADDR(1)",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(1),
        SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(1),
        HoldLow        => thold_RADDR_RCLK_posedge_posedge(1),
        HoldHigh       => thold_RADDR_RCLK_negedge_posedge(1),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR2_RCLK_posedge,
        TimingData     => Tmkr_RADDR2_RCLK_posedge,
        TestSignal     => RADDR_ipd(2),
        TestSignalName => "RADDR(2)",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(2),
        SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(2),
        HoldLow        => thold_RADDR_RCLK_posedge_posedge(2),
        HoldHigh       => thold_RADDR_RCLK_negedge_posedge(2),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR3_RCLK_posedge,
        TimingData     => Tmkr_RADDR3_RCLK_posedge,
        TestSignal     => RADDR_ipd(3),
        TestSignalName => "RADDR(3)",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(3),
        SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(3),
        HoldLow        => thold_RADDR_RCLK_posedge_posedge(3),
        HoldHigh       => thold_RADDR_RCLK_negedge_posedge(3),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR4_RCLK_posedge,
        TimingData     => Tmkr_RADDR4_RCLK_posedge,
        TestSignal     => RADDR_ipd(4),
        TestSignalName => "RADDR(4)",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(4),
        SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(4),
        HoldLow        => thold_RADDR_RCLK_posedge_posedge(4),
        HoldHigh       => thold_RADDR_RCLK_negedge_posedge(4),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR5_RCLK_posedge,
        TimingData     => Tmkr_RADDR5_RCLK_posedge,
        TestSignal     => RADDR_ipd(5),
        TestSignalName => "RADDR(5)",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(5),
        SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(5),
        HoldLow        => thold_RADDR_RCLK_posedge_posedge(5),
        HoldHigh       => thold_RADDR_RCLK_negedge_posedge(5),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR6_RCLK_posedge,
        TimingData     => Tmkr_RADDR6_RCLK_posedge,
        TestSignal     => RADDR_ipd(6),
        TestSignalName => "RADDR(6)",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(6),
        SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(6),
        HoldLow        => thold_RADDR_RCLK_posedge_posedge(6),
        HoldHigh       => thold_RADDR_RCLK_negedge_posedge(6),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR7_RCLK_posedge,
        TimingData     => Tmkr_RADDR7_RCLK_posedge,
        TestSignal     => RADDR_ipd(7),
        TestSignalName => "RADDR(7)",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(7),
        SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(7),
        HoldLow        => thold_RADDR_RCLK_posedge_posedge(7),
        HoldHigh       => thold_RADDR_RCLK_negedge_posedge(7),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_RCLKE_RCLK_posedge,
        TimingData     => Tmkr_RCLKE_RCLK_posedge,
        TestSignal     => RCLKE_ipd,
        TestSignalName => "RCLKE",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RCLKE_RCLK_posedge_posedge,
        SetupLow       => tsetup_RCLKE_RCLK_negedge_posedge,
        HoldLow        => thold_RCLKE_RCLK_posedge_posedge,
        HoldHigh       => thold_RCLKE_RCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_RE_RCLK_posedge,
        TimingData     => Tmkr_RE_RCLK_posedge,
        TestSignal     => RCLK_ipd,
        TestSignalName => "RCLK",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RE_RCLK_posedge_posedge,
        SetupLow       => tsetup_RE_RCLK_negedge_posedge,
        HoldLow        => thold_RE_RCLK_posedge_posedge,
        HoldHigh       => thold_RE_RCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
               

      VitalPeriodPulseCheck (
        Violation      => Pviol_RCLK,
        PeriodData     => PInfo_RCLK,
        TestSignal     => RCLK_ipd,
        TestSignalName => "RCLK",
        TestDelay      => 0 ns,
        Period         => 0 ns,
        PulseWidthHigh => tpw_RCLK_posedge,
        PulseWidthLow  => tpw_RCLK_negedge,
        CheckEnabled   => true,
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);



    end if ;

    Violation  := Pviol_RCLK or
                  Tviol_RADDR0_RCLK_posedge or
                  Tviol_RADDR1_RCLK_posedge or
                  Tviol_RADDR2_RCLK_posedge or
                  Tviol_RADDR3_RCLK_posedge or
                  Tviol_RADDR4_RCLK_posedge or
                  Tviol_RADDR5_RCLK_posedge or
                  Tviol_RADDR6_RCLK_posedge or
                  Tviol_RADDR7_RCLK_posedge or
                  Tviol_RCLKE_RCLK_posedge or
                  Tviol_RE_RCLK_posedge;

    RDATA_zd(0) := Violation xor RDATA_zd(0) ;
    RDATA_zd(1) := Violation xor RDATA_zd(1) ;
    RDATA_zd(2) := Violation xor RDATA_zd(2) ;
    RDATA_zd(3) := Violation xor RDATA_zd(3) ;
    RDATA_zd(4) := Violation xor RDATA_zd(4) ;
    RDATA_zd(5) := Violation xor RDATA_zd(5) ;
    RDATA_zd(6) := Violation xor RDATA_zd(6) ;
    RDATA_zd(7) := Violation xor RDATA_zd(7) ;
    RDATA_zd(8) := Violation xor RDATA_zd(8) ;
    RDATA_zd(9) := Violation xor RDATA_zd(9) ;
    RDATA_zd(10) := Violation xor RDATA_zd(10) ;
    RDATA_zd(11) := Violation xor RDATA_zd(11) ;
    RDATA_zd(12) := Violation xor RDATA_zd(12) ;
    RDATA_zd(13) := Violation xor RDATA_zd(13) ;
    RDATA_zd(14) := Violation xor RDATA_zd(14) ;
    RDATA_zd(15) := Violation xor RDATA_zd(15) ;
    
    
    
    
    
  ----------------------
  --  Path Delay Section
  ----------------------
    VitalPathDelay01 (
      OutSignal     => RDATA(0),
      GlitchData    => RDATA_GlitchData0,
      OutSignalName => "RDATA(0)",
      OutTemp       => RDATA_zd(0),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(0), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(1),
      GlitchData    => RDATA_GlitchData1,
      OutSignalName => "RDATA(1)",
      OutTemp       => RDATA_zd(1),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(1), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(2),
      GlitchData    => RDATA_GlitchData2,
      OutSignalName => "RDATA(2)",
      OutTemp       => RDATA_zd(2),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(2), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(3),
      GlitchData    => RDATA_GlitchData3,
      OutSignalName => "RDATA(3)",
      OutTemp       => RDATA_zd(3),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(3), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(4),
      GlitchData    => RDATA_GlitchData4,
      OutSignalName => "RDATA(4)",
      OutTemp       => RDATA_zd(4),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(4), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(5),
      GlitchData    => RDATA_GlitchData5,
      OutSignalName => "RDATA(5)",
      OutTemp       => RDATA_zd(5),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(5), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(6),
      GlitchData    => RDATA_GlitchData6,
      OutSignalName => "RDATA(6)",
      OutTemp       => RDATA_zd(6),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(6), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(7),
      GlitchData    => RDATA_GlitchData7,
      OutSignalName => "RDATA(7)",
      OutTemp       => RDATA_zd(7),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(7), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(8),
      GlitchData    => RDATA_GlitchData8,
      OutSignalName => "RDATA(8)",
      OutTemp       => RDATA_zd(8),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(8), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(9),
      GlitchData    => RDATA_GlitchData9,
      OutSignalName => "RDATA(9)",
      OutTemp       => RDATA_zd(9),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(9), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(10),
      GlitchData    => RDATA_GlitchData10,
      OutSignalName => "RDATA(10)",
      OutTemp       => RDATA_zd(10),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(10), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(11),
      GlitchData    => RDATA_GlitchData11,
      OutSignalName => "RDATA(11)",
      OutTemp       => RDATA_zd(11),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(11), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(12),
      GlitchData    => RDATA_GlitchData12,
      OutSignalName => "RDATA(12)",
      OutTemp       => RDATA_zd(12),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(12), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(13),
      GlitchData    => RDATA_GlitchData13,
      OutSignalName => "RDATA(13)",
      OutTemp       => RDATA_zd(13),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(13), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(14),
      GlitchData    => RDATA_GlitchData14,
      OutSignalName => "RDATA(14)",
      OutTemp       => RDATA_zd(14),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(14), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(15),
      GlitchData    => RDATA_GlitchData15,
      OutSignalName => "RDATA(15)",
      OutTemp       => RDATA_zd(15),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(15), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(0),
      GlitchData    => RDATA_GlitchData0,
      OutSignalName => "RDATA(0)",
      OutTemp       => RDATA_zd(0),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(0), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(1),
      GlitchData    => RDATA_GlitchData1,
      OutSignalName => "RDATA(1)",
      OutTemp       => RDATA_zd(1),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(1), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(2),
      GlitchData    => RDATA_GlitchData2,
      OutSignalName => "RDATA(2)",
      OutTemp       => RDATA_zd(2),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(2), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(3),
      GlitchData    => RDATA_GlitchData3,
      OutSignalName => "RDATA(3)",
      OutTemp       => RDATA_zd(3),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(3), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(4),
      GlitchData    => RDATA_GlitchData4,
      OutSignalName => "RDATA(4)",
      OutTemp       => RDATA_zd(4),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(4), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(5),
      GlitchData    => RDATA_GlitchData5,
      OutSignalName => "RDATA(5)",
      OutTemp       => RDATA_zd(5),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(5), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(6),
      GlitchData    => RDATA_GlitchData6,
      OutSignalName => "RDATA(6)",
      OutTemp       => RDATA_zd(6),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(6), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(7),
      GlitchData    => RDATA_GlitchData7,
      OutSignalName => "RDATA(7)",
      OutTemp       => RDATA_zd(7),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(7), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(8),
      GlitchData    => RDATA_GlitchData8,
      OutSignalName => "RDATA(8)",
      OutTemp       => RDATA_zd(8),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(8), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(9),
      GlitchData    => RDATA_GlitchData9,
      OutSignalName => "RDATA(9)",
      OutTemp       => RDATA_zd(9),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(9), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(10),
      GlitchData    => RDATA_GlitchData10,
      OutSignalName => "RDATA(10)",
      OutTemp       => RDATA_zd(10),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(10), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(11),
      GlitchData    => RDATA_GlitchData11,
      OutSignalName => "RDATA(11)",
      OutTemp       => RDATA_zd(11),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(11), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(12),
      GlitchData    => RDATA_GlitchData12,
      OutSignalName => "RDATA(12)",
      OutTemp       => RDATA_zd(12),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(12), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(13),
      GlitchData    => RDATA_GlitchData13,
      OutSignalName => "RDATA(13)",
      OutTemp       => RDATA_zd(13),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(13), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(14),
      GlitchData    => RDATA_GlitchData14,
      OutSignalName => "RDATA(14)",
      OutTemp       => RDATA_zd(14),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(14), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(15),
      GlitchData    => RDATA_GlitchData15,
      OutSignalName => "RDATA(15)",
      OutTemp       => RDATA_zd(15),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(15), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

  end process VITALReadBehavior;



  VITALWriteBehavior : process(WADDR_ipd,WCLK_ipd,WCLKE_ipd,WE_ipd,MASK_ipd) 

       variable Tviol_WADDR0_WCLK_posedge : std_logic := '0';
       variable Tviol_WADDR1_WCLK_posedge : std_logic := '0';
       variable Tviol_WADDR2_WCLK_posedge : std_logic := '0';
       variable Tviol_WADDR3_WCLK_posedge : std_logic := '0';
       variable Tviol_WADDR4_WCLK_posedge : std_logic := '0';
       variable Tviol_WADDR5_WCLK_posedge : std_logic := '0';
       variable Tviol_WADDR6_WCLK_posedge : std_logic := '0';
       variable Tviol_WADDR7_WCLK_posedge : std_logic := '0';
       variable Tviol_WCLKE_WCLK_posedge  : std_logic := '0';
       variable Tviol_WE_WCLK_posedge     : std_logic := '0';
       variable Tviol_WDATA0_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA1_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA2_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA3_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA4_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA5_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA6_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA7_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA8_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA9_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA10_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA11_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA12_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA13_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA14_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA15_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK0_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK1_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK2_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK3_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK4_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK5_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK6_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK7_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK8_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK9_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK10_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK11_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK12_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK13_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK14_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK15_WCLK_posedge : std_logic := '0';


       variable Tmkr_WADDR0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR5_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR6_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR7_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WCLKE_WCLK_posedge  : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WE_WCLK_posedge     : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA5_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA6_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA7_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA8_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA9_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA10_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA11_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA12_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA13_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA14_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA15_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK5_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK6_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK7_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK8_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK9_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK10_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK11_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK12_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK13_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK14_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK15_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;

       variable PViol_WCLK : std_logic := '0';

       variable PInfo_WCLK : VitalPeriodDataType := VitalPeriodDataInit;


       variable Violation     : std_logic  := '0';

       variable MEM_temp : std_logic_vector(4095 downto 0) := To_StdLogicVector(INIT_F) &
                                                              To_StdLogicVector(INIT_E) &
                                                              To_StdLogicVector(INIT_D) &
                                                              To_StdLogicVector(INIT_C) &
                                                              To_StdLogicVector(INIT_B) &
                                                              To_StdLogicVector(INIT_A) &
                                                              To_StdLogicVector(INIT_9) &
                                                              To_StdLogicVector(INIT_8) &
                                                              To_StdLogicVector(INIT_7) &
                                                              To_StdLogicVector(INIT_6) &
                                                              To_StdLogicVector(INIT_5) &
                                                              To_StdLogicVector(INIT_4) &
                                                              To_StdLogicVector(INIT_3) &
                                                              To_StdLogicVector(INIT_2) &
                                                              To_StdLogicVector(INIT_1) &
                                                              To_StdLogicVector(INIT_0);
       
  begin

    Violation  := Pviol_WCLK or
                  Tviol_WADDR0_WCLK_posedge or
                  Tviol_WADDR1_WCLK_posedge or
                  Tviol_WADDR2_WCLK_posedge or
                  Tviol_WADDR3_WCLK_posedge or
                  Tviol_WADDR4_WCLK_posedge or
                  Tviol_WADDR5_WCLK_posedge or
                  Tviol_WADDR6_WCLK_posedge or
                  Tviol_WADDR7_WCLK_posedge or
                  Tviol_WCLKE_WCLK_posedge or
                  Tviol_WE_WCLK_posedge or
                  Tviol_WDATA0_WCLK_posedge or
                  Tviol_WDATA1_WCLK_posedge or
                  Tviol_WDATA2_WCLK_posedge or
                  Tviol_WDATA3_WCLK_posedge or
                  Tviol_WDATA4_WCLK_posedge or
                  Tviol_WDATA5_WCLK_posedge or
                  Tviol_WDATA6_WCLK_posedge or
                  Tviol_WDATA7_WCLK_posedge or
                  Tviol_WDATA8_WCLK_posedge or
                  Tviol_WDATA9_WCLK_posedge or
                  Tviol_WDATA10_WCLK_posedge or
                  Tviol_WDATA11_WCLK_posedge or
                  Tviol_WDATA12_WCLK_posedge or
                  Tviol_WDATA13_WCLK_posedge or
                  Tviol_WDATA14_WCLK_posedge or
                  Tviol_WDATA15_WCLK_posedge or
                  Tviol_MASK0_WCLK_posedge or
                  Tviol_MASK1_WCLK_posedge or
                  Tviol_MASK2_WCLK_posedge or
                  Tviol_MASK3_WCLK_posedge or
                  Tviol_MASK4_WCLK_posedge or
                  Tviol_MASK5_WCLK_posedge or
                  Tviol_MASK6_WCLK_posedge or
                  Tviol_MASK7_WCLK_posedge or
                  Tviol_MASK8_WCLK_posedge or
                  Tviol_MASK9_WCLK_posedge or
                  Tviol_MASK10_WCLK_posedge or
                  Tviol_MASK11_WCLK_posedge or
                  Tviol_MASK12_WCLK_posedge or
                  Tviol_MASK13_WCLK_posedge or
                  Tviol_MASK14_WCLK_posedge or
                  Tviol_MASK15_WCLK_posedge;
 
-------------------------
--  Functionality Section
-------------------------

    WADDR_in <= conv_integer(WADDR_ipd) ;
  
    if (Violation = '1') then
       MEM <= (others => 'X') ;
    elsif ( WCLK_ipd'event and (WCLK_ipd = '1') and (WCLKE_ipd = '1' or WCLKE_ipd = 'H') and (WE_ipd = '1') ) then
       for i in 0 to 15 loop
         if (MASK_ipd(i) = '0') then           
            MEM_temp(16*WADDR_in + i ) := WDATA_ipd(i) ;
         end if ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;

------------------------
--  Timing Check Section
------------------------
    if (TimingChecksOn) then
      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR0_WCLK_posedge,
        TimingData     => Tmkr_WADDR0_WCLK_posedge,
        TestSignal     => WADDR_ipd(0),
        TestSignalName => "WADDR(0)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(0),
        SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(0),
        HoldLow        => thold_WADDR_WCLK_posedge_posedge(0),
        HoldHigh       => thold_WADDR_WCLK_negedge_posedge(0),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR1_WCLK_posedge,
        TimingData     => Tmkr_WADDR1_WCLK_posedge,
        TestSignal     => WADDR_ipd(1),
        TestSignalName => "WADDR(1)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(1),
        SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(1),
        HoldLow        => thold_WADDR_WCLK_posedge_posedge(1),
        HoldHigh       => thold_WADDR_WCLK_negedge_posedge(1),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR2_WCLK_posedge,
        TimingData     => Tmkr_WADDR2_WCLK_posedge,
        TestSignal     => WADDR_ipd(2),
        TestSignalName => "WADDR(2)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(2),
        SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(2),
        HoldLow        => thold_WADDR_WCLK_posedge_posedge(2),
        HoldHigh       => thold_WADDR_WCLK_negedge_posedge(2),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR3_WCLK_posedge,
        TimingData     => Tmkr_WADDR3_WCLK_posedge,
        TestSignal     => WADDR_ipd(3),
        TestSignalName => "WADDR(3)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(3),
        SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(3),
        HoldLow        => thold_WADDR_WCLK_posedge_posedge(3),
        HoldHigh       => thold_WADDR_WCLK_negedge_posedge(3),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR4_WCLK_posedge,
        TimingData     => Tmkr_WADDR4_WCLK_posedge,
        TestSignal     => WADDR_ipd(4),
        TestSignalName => "WADDR(4)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(4),
        SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(4),
        HoldLow        => thold_WADDR_WCLK_posedge_posedge(4),
        HoldHigh       => thold_WADDR_WCLK_negedge_posedge(4),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR5_WCLK_posedge,
        TimingData     => Tmkr_WADDR5_WCLK_posedge,
        TestSignal     => WADDR_ipd(5),
        TestSignalName => "WADDR(5)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(5),
        SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(5),
        HoldLow        => thold_WADDR_WCLK_posedge_posedge(5),
        HoldHigh       => thold_WADDR_WCLK_negedge_posedge(5),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR6_WCLK_posedge,
        TimingData     => Tmkr_WADDR6_WCLK_posedge,
        TestSignal     => WADDR_ipd(6),
        TestSignalName => "WADDR(6)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(6),
        SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(6),
        HoldLow        => thold_WADDR_WCLK_posedge_posedge(6),
        HoldHigh       => thold_WADDR_WCLK_negedge_posedge(6),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR7_WCLK_posedge,
        TimingData     => Tmkr_WADDR7_WCLK_posedge,
        TestSignal     => WADDR_ipd(7),
        TestSignalName => "WADDR(7)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(7),
        SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(7),
        HoldLow        => thold_WADDR_WCLK_posedge_posedge(7),
        HoldHigh       => thold_WADDR_WCLK_negedge_posedge(7),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WCLKE_WCLK_posedge,
        TimingData     => Tmkr_WCLKE_WCLK_posedge,
        TestSignal     => WCLKE_ipd,
        TestSignalName => "WCLKE",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WCLKE_WCLK_posedge_posedge,
        SetupLow       => tsetup_WCLKE_WCLK_negedge_posedge,
        HoldLow        => thold_WCLKE_WCLK_posedge_posedge,
        HoldHigh       => thold_WCLKE_WCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WE_WCLK_posedge,
        TimingData     => Tmkr_WE_WCLK_posedge,
        TestSignal     => WCLK_ipd,
        TestSignalName => "WCLK",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WE_WCLK_posedge_posedge,
        SetupLow       => tsetup_WE_WCLK_negedge_posedge,
        HoldLow        => thold_WE_WCLK_posedge_posedge,
        HoldHigh       => thold_WE_WCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
       VitalSetupHoldCheck (
        Violation      => Tviol_WDATA0_WCLK_posedge,
        TimingData     => Tmkr_WDATA0_WCLK_posedge,
        TestSignal     => WDATA_ipd(0),
        TestSignalName => "WDATA(0)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(0),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(0),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(0),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(0),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA1_WCLK_posedge,
        TimingData     => Tmkr_WDATA1_WCLK_posedge,
        TestSignal     => WDATA_ipd(1),
        TestSignalName => "WDATA(1)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(1),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(1),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(1),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(1),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA2_WCLK_posedge,
        TimingData     => Tmkr_WDATA2_WCLK_posedge,
        TestSignal     => WDATA_ipd(2),
        TestSignalName => "WDATA(2)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(2),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(2),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(2),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(2),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA3_WCLK_posedge,
        TimingData     => Tmkr_WDATA3_WCLK_posedge,
        TestSignal     => WDATA_ipd(3),
        TestSignalName => "WDATA(3)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(3),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(3),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(3),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(3),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA4_WCLK_posedge,
        TimingData     => Tmkr_WDATA4_WCLK_posedge,
        TestSignal     => WDATA_ipd(4),
        TestSignalName => "WDATA(4)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(4),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(4),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(4),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(4),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA5_WCLK_posedge,
        TimingData     => Tmkr_WDATA5_WCLK_posedge,
        TestSignal     => WDATA_ipd(5),
        TestSignalName => "WDATA(5)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(5),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(5),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(5),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(5),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA6_WCLK_posedge,
        TimingData     => Tmkr_WDATA6_WCLK_posedge,
        TestSignal     => WDATA_ipd(6),
        TestSignalName => "WDATA(6)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(6),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(6),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(6),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(6),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA7_WCLK_posedge,
        TimingData     => Tmkr_WDATA7_WCLK_posedge,
        TestSignal     => WDATA_ipd(7),
        TestSignalName => "WDATA(7)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(7),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(7),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(7),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(7),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

       VitalSetupHoldCheck (
        Violation      => Tviol_WDATA8_WCLK_posedge,
        TimingData     => Tmkr_WDATA8_WCLK_posedge,
        TestSignal     => WDATA_ipd(8),
        TestSignalName => "WDATA(8)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(8),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(8),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(8),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(8),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA9_WCLK_posedge,
        TimingData     => Tmkr_WDATA9_WCLK_posedge,
        TestSignal     => WDATA_ipd(9),
        TestSignalName => "WDATA(9)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(9),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(9),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(9),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(9),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA10_WCLK_posedge,
        TimingData     => Tmkr_WDATA10_WCLK_posedge,
        TestSignal     => WDATA_ipd(10),
        TestSignalName => "WDATA(10)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(10),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(10),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(10),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(10),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA11_WCLK_posedge,
        TimingData     => Tmkr_WDATA11_WCLK_posedge,
        TestSignal     => WDATA_ipd(11),
        TestSignalName => "WDATA(11)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(11),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(11),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(11),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(11),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA12_WCLK_posedge,
        TimingData     => Tmkr_WDATA12_WCLK_posedge,
        TestSignal     => WDATA_ipd(12),
        TestSignalName => "WDATA(12)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(12),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(12),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(12),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(12),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA13_WCLK_posedge,
        TimingData     => Tmkr_WDATA13_WCLK_posedge,
        TestSignal     => WDATA_ipd(13),
        TestSignalName => "WDATA(13)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(13),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(13),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(13),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(13),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA14_WCLK_posedge,
        TimingData     => Tmkr_WDATA14_WCLK_posedge,
        TestSignal     => WDATA_ipd(14),
        TestSignalName => "WDATA(14)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(14),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(14),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(14),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(14),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA15_WCLK_posedge,
        TimingData     => Tmkr_WDATA15_WCLK_posedge,
        TestSignal     => WDATA_ipd(15),
        TestSignalName => "WDATA(15)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(15),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(15),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(15),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(15),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

       VitalSetupHoldCheck (
        Violation      => Tviol_MASK0_WCLK_posedge,
        TimingData     => Tmkr_MASK0_WCLK_posedge,
        TestSignal     => MASK_ipd(0),
        TestSignalName => "MASK(0)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(0),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(0),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(0),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(0),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK1_WCLK_posedge,
        TimingData     => Tmkr_MASK1_WCLK_posedge,
        TestSignal     => MASK_ipd(1),
        TestSignalName => "MASK(1)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(1),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(1),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(1),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(1),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK2_WCLK_posedge,
        TimingData     => Tmkr_MASK2_WCLK_posedge,
        TestSignal     => MASK_ipd(2),
        TestSignalName => "MASK(2)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(2),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(2),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(2),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(2),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK3_WCLK_posedge,
        TimingData     => Tmkr_MASK3_WCLK_posedge,
        TestSignal     => MASK_ipd(3),
        TestSignalName => "MASK(3)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(3),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(3),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(3),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(3),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK4_WCLK_posedge,
        TimingData     => Tmkr_MASK4_WCLK_posedge,
        TestSignal     => MASK_ipd(4),
        TestSignalName => "MASK(4)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(4),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(4),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(4),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(4),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_MASK5_WCLK_posedge,
        TimingData     => Tmkr_MASK5_WCLK_posedge,
        TestSignal     => MASK_ipd(5),
        TestSignalName => "MASK(5)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(5),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(5),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(5),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(5),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_MASK6_WCLK_posedge,
        TimingData     => Tmkr_MASK6_WCLK_posedge,
        TestSignal     => MASK_ipd(6),
        TestSignalName => "MASK(6)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(6),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(6),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(6),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(6),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_MASK7_WCLK_posedge,
        TimingData     => Tmkr_MASK7_WCLK_posedge,
        TestSignal     => MASK_ipd(7),
        TestSignalName => "MASK(7)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(7),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(7),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(7),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(7),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

       VitalSetupHoldCheck (
        Violation      => Tviol_MASK8_WCLK_posedge,
        TimingData     => Tmkr_MASK8_WCLK_posedge,
        TestSignal     => MASK_ipd(8),
        TestSignalName => "MASK(8)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(8),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(8),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(8),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(8),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK9_WCLK_posedge,
        TimingData     => Tmkr_MASK9_WCLK_posedge,
        TestSignal     => MASK_ipd(9),
        TestSignalName => "MASK(9)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(9),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(9),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(9),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(9),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK10_WCLK_posedge,
        TimingData     => Tmkr_MASK10_WCLK_posedge,
        TestSignal     => MASK_ipd(10),
        TestSignalName => "MASK(10)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(10),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(10),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(10),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(10),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK11_WCLK_posedge,
        TimingData     => Tmkr_MASK11_WCLK_posedge,
        TestSignal     => MASK_ipd(11),
        TestSignalName => "MASK(11)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(11),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(11),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(11),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(11),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK12_WCLK_posedge,
        TimingData     => Tmkr_MASK12_WCLK_posedge,
        TestSignal     => MASK_ipd(12),
        TestSignalName => "MASK(12)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(12),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(12),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(12),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(12),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_MASK13_WCLK_posedge,
        TimingData     => Tmkr_MASK13_WCLK_posedge,
        TestSignal     => MASK_ipd(13),
        TestSignalName => "MASK(13)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(13),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(13),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(13),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(13),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_MASK14_WCLK_posedge,
        TimingData     => Tmkr_MASK14_WCLK_posedge,
        TestSignal     => MASK_ipd(14),
        TestSignalName => "MASK(14)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(14),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(14),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(14),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(14),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_MASK15_WCLK_posedge,
        TimingData     => Tmkr_MASK15_WCLK_posedge,
        TestSignal     => MASK_ipd(15),
        TestSignalName => "MASK(15)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(15),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(15),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(15),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(15),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
   

      VitalPeriodPulseCheck (
        Violation      => Pviol_WCLK,
        PeriodData     => PInfo_WCLK,
        TestSignal     => WCLK_ipd,
        TestSignalName => "WCLK",
        TestDelay      => 0 ns,
        Period         => 0 ns,
        PulseWidthHigh => tpw_WCLK_posedge,
        PulseWidthLow  => tpw_WCLK_negedge,
        CheckEnabled   => true,
        HeaderMsg      => "/SB_RAM4K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);



    end if ;

  end process VITALWriteBehavior;

end SB_RAM4K_V;

--///////////////////////////////////// ---
	--- ICE40 RAM Primitives ---
--///////////////////////////////////// ---


---------------------------------------
	--- SB_RAM256x16
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM256x16 is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 15  downto 0) ;
                RCLK  : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'L';
                RADDR : in  std_logic_vector( 7  downto 0) ;
                WCLK  : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'L';
                WADDR : in  std_logic_vector( 7  downto 0) ;
                MASK  : in  std_logic_vector( 15  downto 0) ;
                WDATA : in  std_logic_vector( 15  downto 0)
               );
  
  
end SB_RAM256x16;

architecture SB_RAM256x16_ARCH of SB_RAM256x16 is

  signal MEM : std_logic_vector(4095 downto 0) ;


  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLK)
  variable WADDR_in : integer range 0 to 255 ;

    variable MEM_temp : std_logic_vector(4095 downto 0) := To_StdLogicVector(INIT_F) &
                                                  To_StdLogicVector(INIT_E) &
                                                  To_StdLogicVector(INIT_D) &
                                                  To_StdLogicVector(INIT_C) &
                                                  To_StdLogicVector(INIT_B) &
                                                  To_StdLogicVector(INIT_A) &
                                                  To_StdLogicVector(INIT_9) &
                                                  To_StdLogicVector(INIT_8) &
                                                  To_StdLogicVector(INIT_7) &
                                                  To_StdLogicVector(INIT_6) &
                                                  To_StdLogicVector(INIT_5) &
                                                  To_StdLogicVector(INIT_4) &
                                                  To_StdLogicVector(INIT_3) &
                                                  To_StdLogicVector(INIT_2) &
                                                  To_StdLogicVector(INIT_1) &
                                                  To_StdLogicVector(INIT_0) ;

  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLK'event and (WCLK = '1') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 15 loop
         if (MASK(i) = '0') then
            MEM_temp(16*WADDR_in + i )  := WDATA(i) ;
         end if ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;


  end process ;


  ReadBehavior : process(RCLK)
  
    variable RADDR_in : integer range 0 to 255 ;
    variable RDATA_temp : std_logic_vector( 15  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLK'event and (RCLK = '1') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 15 loop
            RDATA_temp(i ) := MEM(16*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;


  end process ;
end SB_RAM256x16_ARCH;   --- SB_RAM256x16


---------------------------------------
	--- SB_RAM256x16NR
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM256x16NR is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 15  downto 0) ;
                RCLKN : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'L';
                RADDR : in  std_logic_vector( 7  downto 0) ;
                WCLK  : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'L';
                WADDR : in  std_logic_vector( 7  downto 0) ;
                MASK  : in  std_logic_vector( 15  downto 0) ;
                WDATA : in  std_logic_vector( 15  downto 0)
               );
  
  
end SB_RAM256x16NR;

architecture SB_RAM256x16NR_ARCH of SB_RAM256x16NR is
  signal MEM : std_logic_vector(4095 downto 0) ;


  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLK)
  variable WADDR_in : integer range 0 to 255 ;

    variable MEM_temp : std_logic_vector(4095 downto 0) := To_StdLogicVector(INIT_F) &
                                                  To_StdLogicVector(INIT_E) &
                                                  To_StdLogicVector(INIT_D) &
                                                  To_StdLogicVector(INIT_C) &
                                                  To_StdLogicVector(INIT_B) &
                                                  To_StdLogicVector(INIT_A) &
                                                  To_StdLogicVector(INIT_9) &
                                                  To_StdLogicVector(INIT_8) &
                                                  To_StdLogicVector(INIT_7) &
                                                  To_StdLogicVector(INIT_6) &
                                                  To_StdLogicVector(INIT_5) &
                                                  To_StdLogicVector(INIT_4) &
                                                  To_StdLogicVector(INIT_3) &
                                                  To_StdLogicVector(INIT_2) &
                                                  To_StdLogicVector(INIT_1) &
                                                  To_StdLogicVector(INIT_0) ;

  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLK'event and (WCLK = '1') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 15 loop
         if (MASK(i) = '0') then
            MEM_temp(16*WADDR_in + i )  := WDATA(i) ;
         end if ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;


  end process ;


  ReadBehavior : process(RCLKN)
  
    variable RADDR_in : integer range 0 to 255 ;
    variable RDATA_temp : std_logic_vector( 15  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLKN'event and (RCLKN = '0') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 15 loop
            RDATA_temp(i ) := MEM(16*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;


  end process ;
end SB_RAM256x16NR_ARCH;   --- SB_RAM256x16NR


---------------------------------------
	--- SB_RAM256x16NW
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM256x16NW is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 15  downto 0) ;
                RCLK  : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'L';
                RADDR : in  std_logic_vector( 7  downto 0) ;
                WCLKN : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'L';
                WADDR : in  std_logic_vector( 7  downto 0) ;
                MASK  : in  std_logic_vector( 15  downto 0) ;
                WDATA : in  std_logic_vector( 15  downto 0)
               );
  
  
end SB_RAM256X16NW;

architecture SB_RAM256x16NW_ARCH of SB_RAM256x16NW is
  signal MEM : std_logic_vector(4095 downto 0) ;


  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLKN)
  variable WADDR_in : integer range 0 to 255 ;

    variable MEM_temp : std_logic_vector(4095 downto 0) := To_StdLogicVector(INIT_F) &
                                                  To_StdLogicVector(INIT_E) &
                                                  To_StdLogicVector(INIT_D) &
                                                  To_StdLogicVector(INIT_C) &
                                                  To_StdLogicVector(INIT_B) &
                                                  To_StdLogicVector(INIT_A) &
                                                  To_StdLogicVector(INIT_9) &
                                                  To_StdLogicVector(INIT_8) &
                                                  To_StdLogicVector(INIT_7) &
                                                  To_StdLogicVector(INIT_6) &
                                                  To_StdLogicVector(INIT_5) &
                                                  To_StdLogicVector(INIT_4) &
                                                  To_StdLogicVector(INIT_3) &
                                                  To_StdLogicVector(INIT_2) &
                                                  To_StdLogicVector(INIT_1) &
                                                  To_StdLogicVector(INIT_0) ;

  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLKN'event and (WCLKN = '0') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 15 loop
         if (MASK(i) = '0') then
            MEM_temp(16*WADDR_in + i )  := WDATA(i) ;
         end if ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;


  end process ;


  ReadBehavior : process(RCLK)
  
    variable RADDR_in : integer range 0 to 255 ;
    variable RDATA_temp : std_logic_vector( 15  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLK'event and (RCLK = '1') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 15 loop
            RDATA_temp(i ) := MEM(16*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;
    end process;

end SB_RAM256x16NW_ARCH;   --- SB_RAM256x16NW



---------------------------------------
	--- SB_RAM256x16NRNW
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM256x16NRNW is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 15  downto 0) ;
                RCLKN : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'L';
                RADDR : in  std_logic_vector( 7  downto 0) ;
                WCLKN : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'L';
                WADDR : in  std_logic_vector( 7  downto 0) ;
                MASK  : in  std_logic_vector( 15  downto 0) ;
                WDATA : in  std_logic_vector( 15  downto 0)
               );
  
  
end SB_RAM256x16NRNW;

architecture SB_RAM256x16NRNW_ARCH of SB_RAM256x16NRNW is
  signal MEM : std_logic_vector(4095 downto 0) ;


  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLKN)
  variable WADDR_in : integer range 0 to 255 ;

    variable MEM_temp : std_logic_vector(4095 downto 0) := To_StdLogicVector(INIT_F) &
                                                  To_StdLogicVector(INIT_E) &
                                                  To_StdLogicVector(INIT_D) &
                                                  To_StdLogicVector(INIT_C) &
                                                  To_StdLogicVector(INIT_B) &
                                                  To_StdLogicVector(INIT_A) &
                                                  To_StdLogicVector(INIT_9) &
                                                  To_StdLogicVector(INIT_8) &
                                                  To_StdLogicVector(INIT_7) &
                                                  To_StdLogicVector(INIT_6) &
                                                  To_StdLogicVector(INIT_5) &
                                                  To_StdLogicVector(INIT_4) &
                                                  To_StdLogicVector(INIT_3) &
                                                  To_StdLogicVector(INIT_2) &
                                                  To_StdLogicVector(INIT_1) &
                                                  To_StdLogicVector(INIT_0) ;

  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLKN'event and (WCLKN = '0') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 15 loop
         if (MASK(i) = '0') then
            MEM_temp(16*WADDR_in + i )  := WDATA(i) ;
         end if ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;


  end process ;


  ReadBehavior : process(RCLKN)
  
    variable RADDR_in : integer range 0 to 255 ;
    variable RDATA_temp : std_logic_vector( 15  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLKN'event and (RCLKN = '0') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 15 loop
            RDATA_temp(i ) := MEM(16*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;


  end process ;
end SB_RAM256x16NRNW_ARCH;   --- SB_RAM256x16NRNW


---------------------------------------
	--- SB_RAM512x8
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM512x8 is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 7  downto 0) ;
                RCLK  : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'L';
                RADDR : in  std_logic_vector( 8  downto 0) ;
                WCLK  : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'L';
                WADDR : in  std_logic_vector( 8  downto 0) ;
                WDATA : in  std_logic_vector( 7  downto 0)
               );
  
  
end SB_RAM512x8;

architecture SB_RAM512x8_ARCH of SB_RAM512x8 is

  signal MEM : std_logic_vector(4095 downto 0) ;


  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLK)

  variable WADDR_in : integer range 0 to 511 ;
    variable MEM_temp : std_logic_vector(4095 downto 0) := To_StdLogicVector(INIT_F) &
                                                  To_StdLogicVector(INIT_E) &
                                                  To_StdLogicVector(INIT_D) &
                                                  To_StdLogicVector(INIT_C) &
                                                  To_StdLogicVector(INIT_B) &
                                                  To_StdLogicVector(INIT_A) &
                                                  To_StdLogicVector(INIT_9) &
                                                  To_StdLogicVector(INIT_8) &
                                                  To_StdLogicVector(INIT_7) &
                                                  To_StdLogicVector(INIT_6) &
                                                  To_StdLogicVector(INIT_5) &
                                                  To_StdLogicVector(INIT_4) &
                                                  To_StdLogicVector(INIT_3) &
                                                  To_StdLogicVector(INIT_2) &
                                                  To_StdLogicVector(INIT_1) &
                                                  To_StdLogicVector(INIT_0) ;

  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLK'event and (WCLK = '1') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 7 loop
            MEM_temp(8*WADDR_in + i )  := WDATA(i) ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;


  end process ;


  ReadBehavior : process(RCLK)
  
   variable RADDR_in : integer range 0 to 511 ;
    variable RDATA_temp : std_logic_vector( 7  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLK'event and (RCLK = '1') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 7 loop
            RDATA_temp(i ) := MEM(8*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;


  end process ;
end SB_RAM512x8_ARCH;   --- SB_RAM512x8



---------------------------------------
	--- SB_RAM512x8NR
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM512x8NR is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 7  downto 0) ;
                RCLKN : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'L';
                RADDR : in  std_logic_vector( 8  downto 0) ;
                WCLK  : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'L';
                WADDR : in  std_logic_vector( 8  downto 0) ;
                WDATA : in  std_logic_vector( 7  downto 0)
               );
  
  
end SB_RAM512x8NR;

architecture SB_RAM512x8NR_ARCH of SB_RAM512x8NR is

  signal MEM : std_logic_vector(4095 downto 0) ;


  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLK)

  variable WADDR_in : integer range 0 to 511 ;
    variable MEM_temp : std_logic_vector(4095 downto 0) := To_StdLogicVector(INIT_F) &
                                                  To_StdLogicVector(INIT_E) &
                                                  To_StdLogicVector(INIT_D) &
                                                  To_StdLogicVector(INIT_C) &
                                                  To_StdLogicVector(INIT_B) &
                                                  To_StdLogicVector(INIT_A) &
                                                  To_StdLogicVector(INIT_9) &
                                                  To_StdLogicVector(INIT_8) &
                                                  To_StdLogicVector(INIT_7) &
                                                  To_StdLogicVector(INIT_6) &
                                                  To_StdLogicVector(INIT_5) &
                                                  To_StdLogicVector(INIT_4) &
                                                  To_StdLogicVector(INIT_3) &
                                                  To_StdLogicVector(INIT_2) &
                                                  To_StdLogicVector(INIT_1) &
                                                  To_StdLogicVector(INIT_0) ;

  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLK'event and (WCLK = '1') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 7 loop
            MEM_temp(8*WADDR_in + i )  := WDATA(i) ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;


  end process ;


  ReadBehavior : process(RCLKN)
  
    variable RADDR_in : integer range 0 to 511 ;
    variable RDATA_temp : std_logic_vector( 7  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLKN'event and (RCLKN = '0') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 7 loop
            RDATA_temp(i ) := MEM(8*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;


  end process ;
end SB_RAM512x8NR_ARCH;   --- SB_RAM512x8NR



---------------------------------------
	--- SB_RAM512x8NW
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM512x8NW is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 7  downto 0) ;
                RCLK  : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'L';
                RADDR : in  std_logic_vector( 8  downto 0) ;
                WCLKN : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'L';
                WADDR : in  std_logic_vector( 8  downto 0) ;
                WDATA : in  std_logic_vector( 7  downto 0)
               );
  
  
end SB_RAM512x8NW;

architecture SB_RAM512x8NW_ARCH of SB_RAM512x8NW is
  signal MEM : std_logic_vector(4095 downto 0) ;


  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLKN)
  variable WADDR_in : integer range 0 to 511 ;

    variable MEM_temp : std_logic_vector(4095 downto 0) := To_StdLogicVector(INIT_F) &
                                                  To_StdLogicVector(INIT_E) &
                                                  To_StdLogicVector(INIT_D) &
                                                  To_StdLogicVector(INIT_C) &
                                                  To_StdLogicVector(INIT_B) &
                                                  To_StdLogicVector(INIT_A) &
                                                  To_StdLogicVector(INIT_9) &
                                                  To_StdLogicVector(INIT_8) &
                                                  To_StdLogicVector(INIT_7) &
                                                  To_StdLogicVector(INIT_6) &
                                                  To_StdLogicVector(INIT_5) &
                                                  To_StdLogicVector(INIT_4) &
                                                  To_StdLogicVector(INIT_3) &
                                                  To_StdLogicVector(INIT_2) &
                                                  To_StdLogicVector(INIT_1) &
                                                  To_StdLogicVector(INIT_0) ;

  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLKN'event and (WCLKN = '0') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 7 loop
            MEM_temp(8*WADDR_in + i )  := WDATA(i) ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;


  end process ;


  ReadBehavior : process(RCLK)
  
    variable RADDR_in : integer range 0 to 511 ;
    variable RDATA_temp : std_logic_vector( 7  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLK'event and (RCLK = '1') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 7 loop
            RDATA_temp(i ) := MEM(8*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;


  end process ;
end SB_RAM512x8NW_ARCH;   --- SB_RAM512x8NW


---------------------------------------
	--- SB_RAM512x8NRNW
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM512x8NRNW is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 7  downto 0) ;
                RCLKN : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'L';
                RADDR : in  std_logic_vector( 8  downto 0) ;
                WCLKN : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'L';
                WADDR : in  std_logic_vector( 8  downto 0) ;
                WDATA : in  std_logic_vector( 7  downto 0)
               );
  
  
end SB_RAM512x8NRNW;

architecture SB_RAM512x8NRNW_ARCH of SB_RAM512x8NRNW is
  signal MEM : std_logic_vector(4095 downto 0) ;


  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLKN)

  variable WADDR_in : integer range 0 to 511 ;
    variable MEM_temp : std_logic_vector(4095 downto 0) := To_StdLogicVector(INIT_F) &
                                                  To_StdLogicVector(INIT_E) &
                                                  To_StdLogicVector(INIT_D) &
                                                  To_StdLogicVector(INIT_C) &
                                                  To_StdLogicVector(INIT_B) &
                                                  To_StdLogicVector(INIT_A) &
                                                  To_StdLogicVector(INIT_9) &
                                                  To_StdLogicVector(INIT_8) &
                                                  To_StdLogicVector(INIT_7) &
                                                  To_StdLogicVector(INIT_6) &
                                                  To_StdLogicVector(INIT_5) &
                                                  To_StdLogicVector(INIT_4) &
                                                  To_StdLogicVector(INIT_3) &
                                                  To_StdLogicVector(INIT_2) &
                                                  To_StdLogicVector(INIT_1) &
                                                  To_StdLogicVector(INIT_0) ;

  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLKN'event and (WCLKN = '0') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 7 loop
            MEM_temp(8*WADDR_in + i )  := WDATA(i) ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;


  end process ;


  ReadBehavior : process(RCLKN)
  
   variable RADDR_in : integer range 0 to 511 ;
    variable RDATA_temp : std_logic_vector( 7  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLKN'event and (RCLKN = '0') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 7 loop
            RDATA_temp(i ) := MEM(8*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;


  end process ;
end SB_RAM512x8NRNW_ARCH;   --- SB_RAM512x8NRNW


---------------------------------------
	--- SB_RAM1024x4
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM1024x4 is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 3  downto 0) ;
                RCLK  : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'L';
                RADDR : in  std_logic_vector( 9  downto 0) ;
                WCLK  : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'L';
                WADDR : in  std_logic_vector( 9  downto 0) ;
                WDATA : in  std_logic_vector( 3  downto 0)
               );
  
  
end SB_RAM1024x4;

architecture SB_RAM1024x4_ARCH of SB_RAM1024x4 is

  signal MEM : std_logic_vector(4095 downto 0) ;


  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLK)
  variable WADDR_in : integer range 0 to 1023 ;

    variable MEM_temp : std_logic_vector(4095 downto 0) := To_StdLogicVector(INIT_F) &
                                                  To_StdLogicVector(INIT_E) &
                                                  To_StdLogicVector(INIT_D) &
                                                  To_StdLogicVector(INIT_C) &
                                                  To_StdLogicVector(INIT_B) &
                                                  To_StdLogicVector(INIT_A) &
                                                  To_StdLogicVector(INIT_9) &
                                                  To_StdLogicVector(INIT_8) &
                                                  To_StdLogicVector(INIT_7) &
                                                  To_StdLogicVector(INIT_6) &
                                                  To_StdLogicVector(INIT_5) &
                                                  To_StdLogicVector(INIT_4) &
                                                  To_StdLogicVector(INIT_3) &
                                                  To_StdLogicVector(INIT_2) &
                                                  To_StdLogicVector(INIT_1) &
                                                  To_StdLogicVector(INIT_0) ;

  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLK'event and (WCLK = '1') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 3 loop
            MEM_temp(4*WADDR_in + i )  := WDATA(i) ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;


  end process ;


  ReadBehavior : process(RCLK)
  
    variable RADDR_in : integer range 0 to 1023 ;
    variable RDATA_temp : std_logic_vector( 3  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLK'event and (RCLK = '1') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 3 loop
            RDATA_temp(i ) := MEM(4*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;


  end process ;
end SB_RAM1024x4_ARCH;   --- SB_RAM1024x4



---------------------------------------
	--- SB_RAM1024x4NR
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM1024x4NR is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 3  downto 0) ;
                RCLKN : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'L';
                RADDR : in  std_logic_vector( 9  downto 0) ;
                WCLK  : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'L';
                WADDR : in  std_logic_vector( 9  downto 0) ;
                WDATA : in  std_logic_vector( 3  downto 0)
               );
  
  
end SB_RAM1024x4NR;

architecture SB_RAM1024x4NR_ARCH of SB_RAM1024x4NR is
  signal MEM : std_logic_vector(4095 downto 0) ;


  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLK)
  variable WADDR_in : integer range 0 to 1023 ;

    variable MEM_temp : std_logic_vector(4095 downto 0) := To_StdLogicVector(INIT_F) &
                                                  To_StdLogicVector(INIT_E) &
                                                  To_StdLogicVector(INIT_D) &
                                                  To_StdLogicVector(INIT_C) &
                                                  To_StdLogicVector(INIT_B) &
                                                  To_StdLogicVector(INIT_A) &
                                                  To_StdLogicVector(INIT_9) &
                                                  To_StdLogicVector(INIT_8) &
                                                  To_StdLogicVector(INIT_7) &
                                                  To_StdLogicVector(INIT_6) &
                                                  To_StdLogicVector(INIT_5) &
                                                  To_StdLogicVector(INIT_4) &
                                                  To_StdLogicVector(INIT_3) &
                                                  To_StdLogicVector(INIT_2) &
                                                  To_StdLogicVector(INIT_1) &
                                                  To_StdLogicVector(INIT_0) ;

  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLK'event and (WCLK = '1') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 3 loop
            MEM_temp(4*WADDR_in + i )  := WDATA(i) ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;


  end process ;


  ReadBehavior : process(RCLKN)
  
    variable RADDR_in : integer range 0 to 1023 ;
    variable RDATA_temp : std_logic_vector( 3  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLKN'event and (RCLKN = '0') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 3 loop
            RDATA_temp(i ) := MEM(4*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;


  end process ;
end SB_RAM1024x4NR_ARCH;   --- SB_RAM1024x4NR


---------------------------------------
	--- SB_RAM1024x4NW
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM1024x4NW is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 3  downto 0) ;
                RCLK  : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'L';
                RADDR : in  std_logic_vector( 9  downto 0) ;
                WCLKN : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'L';
                WADDR : in  std_logic_vector( 9  downto 0) ;
                WDATA : in  std_logic_vector( 3  downto 0)
               );
  
  
end SB_RAM1024x4NW;

architecture SB_RAM1024x4NW_ARCH of SB_RAM1024x4NW is
  signal MEM : std_logic_vector(4095 downto 0) ;


  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLKN)
  variable WADDR_in : integer range 0 to 1023 ;

    variable MEM_temp : std_logic_vector(4095 downto 0) := To_StdLogicVector(INIT_F) &
                                                  To_StdLogicVector(INIT_E) &
                                                  To_StdLogicVector(INIT_D) &
                                                  To_StdLogicVector(INIT_C) &
                                                  To_StdLogicVector(INIT_B) &
                                                  To_StdLogicVector(INIT_A) &
                                                  To_StdLogicVector(INIT_9) &
                                                  To_StdLogicVector(INIT_8) &
                                                  To_StdLogicVector(INIT_7) &
                                                  To_StdLogicVector(INIT_6) &
                                                  To_StdLogicVector(INIT_5) &
                                                  To_StdLogicVector(INIT_4) &
                                                  To_StdLogicVector(INIT_3) &
                                                  To_StdLogicVector(INIT_2) &
                                                  To_StdLogicVector(INIT_1) &
                                                  To_StdLogicVector(INIT_0) ;

  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLKN'event and (WCLKN = '0') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 3 loop
            MEM_temp(4*WADDR_in + i )  := WDATA(i) ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;


  end process ;


  ReadBehavior : process(RCLK)
  
    variable RADDR_in : integer range 0 to 1023 ;
    variable RDATA_temp : std_logic_vector( 3  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLK'event and (RCLK = '1') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 3 loop
            RDATA_temp(i ) := MEM(4*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;


  end process ;
end SB_RAM1024x4NW_ARCH;   --- SB_RAM1024x4NW


---------------------------------------
	--- SB_RAM1024x4NRNW
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM1024x4NRNW is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 3  downto 0) ;
                RCLKN : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'L';
                RADDR : in  std_logic_vector( 9  downto 0) ;
                WCLKN : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'L';
                WADDR : in  std_logic_vector( 9  downto 0) ;
                WDATA : in  std_logic_vector( 3  downto 0)
               );
  
  
end SB_RAM1024x4NRNW;

architecture SB_RAM1024x4NRNW_ARCH of SB_RAM1024x4NRNW is
  signal MEM : std_logic_vector(4095 downto 0) ;


  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLKN)
  variable WADDR_in : integer range 0 to 1023 ;

    variable MEM_temp : std_logic_vector(4095 downto 0) := To_StdLogicVector(INIT_F) &
                                                  To_StdLogicVector(INIT_E) &
                                                  To_StdLogicVector(INIT_D) &
                                                  To_StdLogicVector(INIT_C) &
                                                  To_StdLogicVector(INIT_B) &
                                                  To_StdLogicVector(INIT_A) &
                                                  To_StdLogicVector(INIT_9) &
                                                  To_StdLogicVector(INIT_8) &
                                                  To_StdLogicVector(INIT_7) &
                                                  To_StdLogicVector(INIT_6) &
                                                  To_StdLogicVector(INIT_5) &
                                                  To_StdLogicVector(INIT_4) &
                                                  To_StdLogicVector(INIT_3) &
                                                  To_StdLogicVector(INIT_2) &
                                                  To_StdLogicVector(INIT_1) &
                                                  To_StdLogicVector(INIT_0) ;

  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLKN'event and (WCLKN = '0') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 3 loop
            MEM_temp(4*WADDR_in + i )  := WDATA(i) ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;


  end process ;


  ReadBehavior : process(RCLKN)
  
    variable RADDR_in : integer range 0 to 1023 ;
    variable RDATA_temp : std_logic_vector( 3  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLKN'event and (RCLKN = '0') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 3 loop
            RDATA_temp(i ) := MEM(4*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;


  end process ;
end SB_RAM1024x4NRNW_ARCH;   --- SB_RAM1024x4NRNW


---------------------------------------
	--- SB_RAM2048x2
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM2048x2 is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 1  downto 0) ;
                RCLK  : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'L';
                RADDR : in  std_logic_vector( 10  downto 0) ;
                WCLK  : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'L';
                WADDR : in  std_logic_vector( 10  downto 0) ;
                WDATA : in  std_logic_vector( 1  downto 0)
               );
  
  
end SB_RAM2048x2;

architecture SB_RAM2048x2_ARCH of SB_RAM2048x2 is

  signal MEM : std_logic_vector(4095 downto 0) ;


  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLK)
  variable WADDR_in : integer range 0 to 2047 ;

    variable MEM_temp : std_logic_vector(4095 downto 0) := To_StdLogicVector(INIT_F) &
                                                  To_StdLogicVector(INIT_E) &
                                                  To_StdLogicVector(INIT_D) &
                                                  To_StdLogicVector(INIT_C) &
                                                  To_StdLogicVector(INIT_B) &
                                                  To_StdLogicVector(INIT_A) &
                                                  To_StdLogicVector(INIT_9) &
                                                  To_StdLogicVector(INIT_8) &
                                                  To_StdLogicVector(INIT_7) &
                                                  To_StdLogicVector(INIT_6) &
                                                  To_StdLogicVector(INIT_5) &
                                                  To_StdLogicVector(INIT_4) &
                                                  To_StdLogicVector(INIT_3) &
                                                  To_StdLogicVector(INIT_2) &
                                                  To_StdLogicVector(INIT_1) &
                                                  To_StdLogicVector(INIT_0) ;

  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLK'event and (WCLK = '1') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 1 loop
            MEM_temp(2*WADDR_in + i )  := WDATA(i) ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;


  end process ;


  ReadBehavior : process(RCLK)
  
    variable RADDR_in : integer range 0 to 2047 ;
    variable RDATA_temp : std_logic_vector( 1  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLK'event and (RCLK = '1') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 1 loop
            RDATA_temp(i ) := MEM(2*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;


  end process ;
end SB_RAM2048x2_ARCH;   --- SB_RAM2048x2


---------------------------------------
	--- SB_RAM2048x2NR
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM2048x2NR is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 1  downto 0) ;
                RCLKN : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'L';
                RADDR : in  std_logic_vector( 10  downto 0) ;
                WCLK  : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'L';
                WADDR : in  std_logic_vector( 10  downto 0) ;
                WDATA : in  std_logic_vector( 1  downto 0)
               );
  
  
end SB_RAM2048x2NR;

architecture SB_RAM2048x2NR_ARCH of SB_RAM2048x2NR is

  signal MEM : std_logic_vector(4095 downto 0) ;


  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLK)
  variable WADDR_in : integer range 0 to 2047 ;

    variable MEM_temp : std_logic_vector(4095 downto 0) := To_StdLogicVector(INIT_F) &
                                                  To_StdLogicVector(INIT_E) &
                                                  To_StdLogicVector(INIT_D) &
                                                  To_StdLogicVector(INIT_C) &
                                                  To_StdLogicVector(INIT_B) &
                                                  To_StdLogicVector(INIT_A) &
                                                  To_StdLogicVector(INIT_9) &
                                                  To_StdLogicVector(INIT_8) &
                                                  To_StdLogicVector(INIT_7) &
                                                  To_StdLogicVector(INIT_6) &
                                                  To_StdLogicVector(INIT_5) &
                                                  To_StdLogicVector(INIT_4) &
                                                  To_StdLogicVector(INIT_3) &
                                                  To_StdLogicVector(INIT_2) &
                                                  To_StdLogicVector(INIT_1) &
                                                  To_StdLogicVector(INIT_0) ;

  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLK'event and (WCLK = '1') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 1 loop
            MEM_temp(2*WADDR_in + i )  := WDATA(i) ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;


  end process ;


  ReadBehavior : process(RCLKN)
  
    variable RADDR_in : integer range 0 to 2047 ;
    variable RDATA_temp : std_logic_vector( 1  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLKN'event and (RCLKN = '0') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 1 loop
            RDATA_temp(i ) := MEM(2*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;


  end process ;
end SB_RAM2048x2NR_ARCH;   --- SB_RAM2048x2NR


---------------------------------------
	--- SB_RAM2048x2NW
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM2048x2NW is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 1  downto 0) ;
                RCLK  : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'L';
                RADDR : in  std_logic_vector( 10  downto 0) ;
                WCLKN : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'L';
                WADDR : in  std_logic_vector( 10  downto 0) ;
                WDATA : in  std_logic_vector( 1  downto 0)
               );
  
  
end SB_RAM2048x2NW;

architecture SB_RAM2048x2NW_ARCH of SB_RAM2048x2NW is

  signal MEM : std_logic_vector(4095 downto 0) ;


  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLKN)
  variable WADDR_in : integer range 0 to 2047 ;

    variable MEM_temp : std_logic_vector(4095 downto 0) := To_StdLogicVector(INIT_F) &
                                                  To_StdLogicVector(INIT_E) &
                                                  To_StdLogicVector(INIT_D) &
                                                  To_StdLogicVector(INIT_C) &
                                                  To_StdLogicVector(INIT_B) &
                                                  To_StdLogicVector(INIT_A) &
                                                  To_StdLogicVector(INIT_9) &
                                                  To_StdLogicVector(INIT_8) &
                                                  To_StdLogicVector(INIT_7) &
                                                  To_StdLogicVector(INIT_6) &
                                                  To_StdLogicVector(INIT_5) &
                                                  To_StdLogicVector(INIT_4) &
                                                  To_StdLogicVector(INIT_3) &
                                                  To_StdLogicVector(INIT_2) &
                                                  To_StdLogicVector(INIT_1) &
                                                  To_StdLogicVector(INIT_0) ;

  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLKN'event and (WCLKN = '0') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 1 loop
            MEM_temp(2*WADDR_in + i )  := WDATA(i) ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;


  end process ;


  ReadBehavior : process(RCLK)
  
    variable RADDR_in : integer range 0 to 2047 ;
    variable RDATA_temp : std_logic_vector( 1  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLK'event and (RCLK = '1') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 1 loop
            RDATA_temp(i ) := MEM(2*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;


  end process ;
end SB_RAM2048x2NW_ARCH;   --- SB_RAM2048x2NW


---------------------------------------
	--- SB_RAM2048x2NRNW
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM2048x2NRNW is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 1  downto 0) ;
                RCLKN : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'L';
                RADDR : in  std_logic_vector( 10  downto 0) ;
                WCLKN : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'L';
                WADDR : in  std_logic_vector( 10  downto 0) ;
                WDATA : in  std_logic_vector( 1  downto 0)
               );
  
  
end SB_RAM2048x2NRNW;

architecture SB_RAM2048x2NRNW_ARCH of SB_RAM2048x2NRNW is

  signal MEM : std_logic_vector(4095 downto 0) ;


  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLKN)
  variable WADDR_in : integer range 0 to 2047 ;

    variable MEM_temp : std_logic_vector(4095 downto 0) := To_StdLogicVector(INIT_F) &
                                                  To_StdLogicVector(INIT_E) &
                                                  To_StdLogicVector(INIT_D) &
                                                  To_StdLogicVector(INIT_C) &
                                                  To_StdLogicVector(INIT_B) &
                                                  To_StdLogicVector(INIT_A) &
                                                  To_StdLogicVector(INIT_9) &
                                                  To_StdLogicVector(INIT_8) &
                                                  To_StdLogicVector(INIT_7) &
                                                  To_StdLogicVector(INIT_6) &
                                                  To_StdLogicVector(INIT_5) &
                                                  To_StdLogicVector(INIT_4) &
                                                  To_StdLogicVector(INIT_3) &
                                                  To_StdLogicVector(INIT_2) &
                                                  To_StdLogicVector(INIT_1) &
                                                  To_StdLogicVector(INIT_0) ;

  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLKN'event and (WCLKN = '0') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 1 loop
            MEM_temp(2*WADDR_in + i )  := WDATA(i) ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;


  end process ;


  ReadBehavior : process(RCLKN)
  
    variable RADDR_in : integer range 0 to 2047 ;
    variable RDATA_temp : std_logic_vector( 1  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLKN'event and (RCLKN = '1') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 1 loop
            RDATA_temp(i ) := MEM(2*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;


  end process ;
end SB_RAM2048x2NRNW_ARCH;   --- SB_RAM2048x2NRNW



---------------------------------------
	--- iCE40P Primitives
---------------------------------------

---------------------------------------
	--- SB_RAM40_4K
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
use IEEE.VITAL_Timing.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM40_4K is

  generic ( 
           TimingChecksOn : boolean := true;
           Xon            : boolean := false;
           MsgOn          : boolean := false;
           
           tipd_RCLK  : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_RCLKE : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_RE    : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_RADDR : VitalDelayArrayType01(10 downto 0) := (others => (0 ns, 0 ns));
           tipd_WCLK  : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_WCLKE : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_WE    : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_WADDR : VitalDelayArrayType01(10 downto 0) := (others => (0 ns, 0 ns));
           tipd_MASK  : VitalDelayArrayType01(15 downto 0) := (others => (0 ns, 0 ns));
           tipd_WDATA : VitalDelayArrayType01(15 downto 0) := (others => (0 ns, 0 ns));
		 		
           tpd_RCLK_RDATA : VitalDelayArrayType01(15 downto 0) := (others => (0 ns, 0 ns));
           tpd_RCLK_RDATA_posedge : VitalDelayArrayType01(15 downto 0) := (others => (0 ns, 0 ns));

           tsetup_RADDR_RCLK_negedge_posedge : VitalDelayArrayType(10 downto 0) := (others => 0 ns);
           tsetup_RADDR_RCLK_posedge_posedge : VitalDelayArrayType(10 downto 0) := (others => 0 ns);
           tsetup_RCLKE_RCLK_negedge_posedge : VitalDelayType                   := 0 ns;
           tsetup_RCLKE_RCLK_posedge_posedge : VitalDelayType                   := 0 ns;
           tsetup_RE_RCLK_negedge_posedge    : VitalDelayType                   := 0 ns;
           tsetup_RE_RCLK_posedge_posedge    : VitalDelayType                   := 0 ns;

           tsetup_WADDR_WCLK_negedge_posedge : VitalDelayArrayType(10 downto 0) := (others => 0 ns);
           tsetup_WADDR_WCLK_posedge_posedge : VitalDelayArrayType(10 downto 0) := (others => 0 ns);
           tsetup_WDATA_WCLK_negedge_posedge : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           tsetup_WDATA_WCLK_posedge_posedge : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           tsetup_WCLKE_WCLK_negedge_posedge : VitalDelayType                   := 0 ns;
           tsetup_WCLKE_WCLK_posedge_posedge : VitalDelayType                   := 0 ns;
           tsetup_WE_WCLK_negedge_posedge    : VitalDelayType                   := 0 ns;
           tsetup_WE_WCLK_posedge_posedge    : VitalDelayType                   := 0 ns;
           tsetup_MASK_WCLK_negedge_posedge  : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           tsetup_MASK_WCLK_posedge_posedge  : VitalDelayArrayType(15 downto 0) := (others => 0 ns);

           thold_RADDR_RCLK_negedge_posedge : VitalDelayArrayType(10 downto 0) := (others => 0 ns);
           thold_RADDR_RCLK_posedge_posedge : VitalDelayArrayType(10 downto 0) := (others => 0 ns);
           thold_RCLKE_RCLK_negedge_posedge : VitalDelayType                   := 0 ns;
           thold_RCLKE_RCLK_posedge_posedge : VitalDelayType                   := 0 ns;
           thold_RE_RCLK_negedge_posedge    : VitalDelayType                   := 0 ns;
           thold_RE_RCLK_posedge_posedge    : VitalDelayType                   := 0 ns;

           thold_WADDR_WCLK_negedge_posedge : VitalDelayArrayType(10 downto 0)  := (others => 0 ns);
           thold_WADDR_WCLK_posedge_posedge : VitalDelayArrayType(10 downto 0)  := (others => 0 ns);
           thold_WDATA_WCLK_negedge_posedge : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           thold_WDATA_WCLK_posedge_posedge : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           thold_WCLKE_WCLK_negedge_posedge : VitalDelayType                   := 0 ns;
           thold_WCLKE_WCLK_posedge_posedge : VitalDelayType                   := 0 ns;
           thold_WE_WCLK_negedge_posedge    : VitalDelayType                   := 0 ns;
           thold_WE_WCLK_posedge_posedge    : VitalDelayType                   := 0 ns;
           thold_MASK_WCLK_negedge_posedge  : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           thold_MASK_WCLK_posedge_posedge  : VitalDelayArrayType(15 downto 0) := (others => 0 ns);

           tpw_RCLK_negedge : VitalDelayType := 0 ns;
           tpw_RCLK_posedge : VitalDelayType := 0 ns;
           tpw_WCLK_negedge : VitalDelayType := 0 ns;
           tpw_WCLK_posedge : VitalDelayType := 0 ns;


  	   WRITE_MODE : integer := 0; -- can be integer 0(256X16 mode) or 1(512X8 mode) or 2(1024X4 mode) or 3(2048X2 mode)
  	   READ_MODE  : integer := 0; -- can be integer 0(256X16 mode) or 1(512X8 mode) or 2(1024X4 mode) or 3(2048X2 mode)
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 15  downto 0) ;
                RCLK  : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'L';
                RADDR : in  std_logic_vector( 10  downto 0) ;
                WCLK  : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'L';
                WADDR : in  std_logic_vector( 10  downto 0) ;
                MASK  : in  std_logic_vector( 15  downto 0) ;
                WDATA : in  std_logic_vector( 15 downto 0)
               );
 
  attribute VITAL_LEVEL0 of SB_RAM40_4K : entity is TRUE;

end SB_RAM40_4K;

architecture SB_RAM40_4K_V of SB_RAM40_4K is

  attribute VITAL_LEVEL0 of SB_RAM40_4K_V  : architecture is TRUE;
  
	 component read_data_decoder 
		generic (
			READ_MODE : integer := 0
		);
		port (
			di	 :  in std_logic_vector (15 downto 0);
			ldo	 :  out std_logic_vector (15 downto 0);
			ai	 :  in std_logic_vector (2 downto 0)
		);
	end component;

	component mask_decoder 
		generic (
			WRITE_MODE : integer := 0 
		);
		port (
			mi	 :  in std_logic_vector (15 downto 0);
			mo	 :  out std_logic_vector (15 downto 0);
			ai	 :  in std_logic_vector (2 downto 0)
		);
	end component;

	component write_data_decoder 
		generic (
			WRITE_MODE  : integer := 0
		);
		port (
			di	 : in std_logic_vector(15 downto 0);
			ldo	 : out std_logic_vector (15 downto 0)
		);
	end component;

	component SB_RAM4K 
		generic (
			INIT_0	   : bit_vector;
			INIT_1	   : bit_vector;
			INIT_2	   : bit_vector;
			INIT_3	   : bit_vector;
			INIT_4	   : bit_vector;
			INIT_5	   : bit_vector;
			INIT_6	   : bit_vector;
			INIT_7	   : bit_vector;
			INIT_8	   : bit_vector;
			INIT_9	   : bit_vector;
			INIT_A	   : bit_vector;
			INIT_B	   : bit_vector;
			INIT_C	   : bit_vector;
			INIT_D	   : bit_vector;
			INIT_E	   : bit_vector;
			INIT_F	   : bit_vector
		);
		port (
			RDATA	   : out std_logic_vector(15 downto 0);
			RCLK	   : in std_logic;
			RCLKE	   : in std_logic;
			RE	   : in std_logic;
			RADDR	   : in std_logic_vector(7 downto 0);
			MASK	   : in std_logic_vector(15 downto 0);
			WDATA	   : in std_logic_vector(15 downto 0);
			WCLK	   : in std_logic;
			WCLKE	   : in std_logic;
			WE	   : in std_logic;
			WADDR	   : in std_logic_vector(7 downto 0)
		);
	end component;


	--- VITAL Signals   
	signal RADDR_ipd : std_logic_vector(10 downto 0)  := (others => 'X');   
	signal RCLK_ipd  : std_logic                    := 'X';
	signal RCLKE_ipd : std_logic                    := 'X';
	signal RE_ipd    : std_logic                    := 'X';

	signal WADDR_ipd : std_logic_vector(10 downto 0)  := (others => 'X');
	signal WCLK_ipd  : std_logic                    := 'X';  
	signal WCLKE_ipd : std_logic                    := 'X';
	signal WE_ipd    : std_logic                    := 'X';
	signal MASK_ipd  : std_logic_vector(15 downto 0) := (others => 'X');
	signal WDATA_ipd : std_logic_vector(15 downto 0) := (others => 'X');

        signal RDATA_zd : std_logic_vector(15 downto 0) := (others => 'X');

	---- Function Signals
	signal RD : std_logic_vector(15 downto 0);
	signal WD : std_logic_vector(15 downto 0);
	signal MASK_RAM : std_logic_vector(15 downto 0);

	signal READ_ADDR_HB : std_logic_vector (2 downto 0);
	signal READ_ADDR_LB : std_logic_vector (7 downto 0);
	signal WRITE_ADDR_LB : std_logic_vector (7 downto 0);
	signal WRITE_ADDR_HB : std_logic_vector (2 downto 0);

	signal READ_ADDR_HB_reg : std_logic_vector (2 downto 0); 
	
begin
	---------------------
	--  Input Wire Delay
	---------------------
	WireDelay : block
	begin
	  RADDR_DELAY : for i in 10 downto 0 generate
	     VitalWireDelay (RADDR_ipd(i), RADDR(i), tipd_RADDR(i));
	  end generate RADDR_DELAY;
	  VitalWireDelay (RCLK_ipd, RCLK, tipd_RCLK);
	  VitalWireDelay (RCLKE_ipd, RCLKE, tipd_RCLKE);
	  VitalWireDelay (RE_ipd, RE, tipd_RE);
	  WADDR_DELAY : for i in 10 downto 0 generate
	     VitalWireDelay (WADDR_ipd(i), WADDR(i), tipd_WADDR(i));
	  end generate WADDR_DELAY;
	  VitalWireDelay (WCLK_ipd, WCLK, tipd_WCLK);
	  VitalWireDelay (WCLKE_ipd, WCLKE, tipd_WCLKE);
	  VitalWireDelay (WE_ipd, WE, tipd_WE);
	  MASK_DELAY : for i in 15 downto 0 generate
	     VitalWireDelay (MASK_ipd(i), MASK(i), tipd_MASK(i));
	  end generate MASK_DELAY;
	  WDATA_DELAY : for i in 15 downto 0 generate
	     VitalWireDelay (WDATA_ipd(i), WDATA(i), tipd_WDATA(i));
	  end generate WDATA_DELAY;
	end block;

	VITALBehavior : block
	begin

	---------------------
	--  Timing Checks
	---------------------
	TimingChecks : process (RADDR_ipd, RCLK_ipd, RCLKE_ipd, RE_ipd, WADDR_ipd, WCLK_ipd, WCLKE_ipd, WE_ipd, MASK_ipd, WDATA_ipd)

	variable Tviol_RADDR0_RCLK_posedge : std_logic := '0';
	variable Tviol_RADDR1_RCLK_posedge : std_logic := '0';
	variable Tviol_RADDR2_RCLK_posedge : std_logic := '0';
	variable Tviol_RADDR3_RCLK_posedge : std_logic := '0';
	variable Tviol_RADDR4_RCLK_posedge : std_logic := '0';
	variable Tviol_RADDR5_RCLK_posedge : std_logic := '0';
	variable Tviol_RADDR6_RCLK_posedge : std_logic := '0';
	variable Tviol_RADDR7_RCLK_posedge : std_logic := '0';
	variable Tviol_RADDR8_RCLK_posedge : std_logic := '0';
	variable Tviol_RADDR9_RCLK_posedge : std_logic := '0';
	variable Tviol_RADDR10_RCLK_posedge : std_logic := '0';
	variable Tviol_RCLKE_RCLK_posedge  : std_logic := '0';
	variable Tviol_RE_RCLK_posedge     : std_logic := '0';

	variable Tmkr_RADDR0_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_RADDR1_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_RADDR2_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_RADDR3_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_RADDR4_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_RADDR5_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_RADDR6_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_RADDR7_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_RADDR8_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_RADDR9_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_RADDR10_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_RCLKE_RCLK_posedge  : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_RE_RCLK_posedge     : VitalTimingDataType := VitalTimingDataInit;

	variable PViol_RCLK : std_logic := '0';

	variable PInfo_RCLK : VitalPeriodDataType ;

        variable Tviol_WADDR0_WCLK_posedge : std_logic := '0';
        variable Tviol_WADDR1_WCLK_posedge : std_logic := '0';
        variable Tviol_WADDR2_WCLK_posedge : std_logic := '0';
        variable Tviol_WADDR3_WCLK_posedge : std_logic := '0';
        variable Tviol_WADDR4_WCLK_posedge : std_logic := '0';
        variable Tviol_WADDR5_WCLK_posedge : std_logic := '0';
        variable Tviol_WADDR6_WCLK_posedge : std_logic := '0';
        variable Tviol_WADDR7_WCLK_posedge : std_logic := '0';
        variable Tviol_WADDR8_WCLK_posedge : std_logic := '0';
        variable Tviol_WADDR9_WCLK_posedge : std_logic := '0';
        variable Tviol_WADDR10_WCLK_posedge : std_logic := '0';
        variable Tviol_WCLKE_WCLK_posedge  : std_logic := '0';
        variable Tviol_WE_WCLK_posedge     : std_logic := '0';
        variable Tviol_WDATA0_WCLK_posedge : std_logic := '0';
        variable Tviol_WDATA1_WCLK_posedge : std_logic := '0';
        variable Tviol_WDATA2_WCLK_posedge : std_logic := '0';
        variable Tviol_WDATA3_WCLK_posedge : std_logic := '0';
        variable Tviol_WDATA4_WCLK_posedge : std_logic := '0';
        variable Tviol_WDATA5_WCLK_posedge : std_logic := '0';
        variable Tviol_WDATA6_WCLK_posedge : std_logic := '0';
        variable Tviol_WDATA7_WCLK_posedge : std_logic := '0';
        variable Tviol_WDATA8_WCLK_posedge : std_logic := '0';
        variable Tviol_WDATA9_WCLK_posedge : std_logic := '0';
        variable Tviol_WDATA10_WCLK_posedge : std_logic := '0';
        variable Tviol_WDATA11_WCLK_posedge : std_logic := '0';
        variable Tviol_WDATA12_WCLK_posedge : std_logic := '0';
        variable Tviol_WDATA13_WCLK_posedge : std_logic := '0';
        variable Tviol_WDATA14_WCLK_posedge : std_logic := '0';
        variable Tviol_WDATA15_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK0_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK1_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK2_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK3_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK4_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK5_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK6_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK7_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK8_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK9_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK10_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK11_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK12_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK13_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK14_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK15_WCLK_posedge : std_logic := '0';


        variable Tmkr_WADDR0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WADDR1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WADDR2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WADDR3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WADDR4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WADDR5_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WADDR6_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WADDR7_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WADDR8_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WADDR9_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WADDR10_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WCLKE_WCLK_posedge  : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WE_WCLK_posedge     : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA5_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA6_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA7_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA8_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA9_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA10_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA11_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA12_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA13_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA14_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA15_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK5_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK6_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK7_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK8_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK9_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK10_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK11_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK12_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK13_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK14_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK15_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;

        variable PViol_WCLK : std_logic := '0';

        variable PInfo_WCLK : VitalPeriodDataType := VitalPeriodDataInit;

	variable Violation     : std_logic  := '0';

	begin

	    if (TimingChecksOn) then
	      VitalSetupHoldCheck (
		Violation      => Tviol_RADDR0_RCLK_posedge,
		TimingData     => Tmkr_RADDR0_RCLK_posedge,
		TestSignal     => RADDR_ipd(0),
		TestSignalName => "RADDR(0)",
		TestDelay      => 0 ns,
		RefSignal      => RCLK_ipd,
		RefSignalName  => "RCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(0),
		SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(0),
		HoldLow        => thold_RADDR_RCLK_posedge_posedge(0),
		HoldHigh       => thold_RADDR_RCLK_negedge_posedge(0),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_RADDR1_RCLK_posedge,
		TimingData     => Tmkr_RADDR1_RCLK_posedge,
		TestSignal     => RADDR_ipd(1),
		TestSignalName => "RADDR(1)",
		TestDelay      => 0 ns,
		RefSignal      => RCLK_ipd,
		RefSignalName  => "RCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(1),
		SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(1),
		HoldLow        => thold_RADDR_RCLK_posedge_posedge(1),
		HoldHigh       => thold_RADDR_RCLK_negedge_posedge(1),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_RADDR2_RCLK_posedge,
		TimingData     => Tmkr_RADDR2_RCLK_posedge,
		TestSignal     => RADDR_ipd(2),
		TestSignalName => "RADDR(2)",
		TestDelay      => 0 ns,
		RefSignal      => RCLK_ipd,
		RefSignalName  => "RCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(2),
		SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(2),
		HoldLow        => thold_RADDR_RCLK_posedge_posedge(2),
		HoldHigh       => thold_RADDR_RCLK_negedge_posedge(2),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_RADDR3_RCLK_posedge,
		TimingData     => Tmkr_RADDR3_RCLK_posedge,
		TestSignal     => RADDR_ipd(3),
		TestSignalName => "RADDR(3)",
		TestDelay      => 0 ns,
		RefSignal      => RCLK_ipd,
		RefSignalName  => "RCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(3),
		SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(3),
		HoldLow        => thold_RADDR_RCLK_posedge_posedge(3),
		HoldHigh       => thold_RADDR_RCLK_negedge_posedge(3),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_RADDR4_RCLK_posedge,
		TimingData     => Tmkr_RADDR4_RCLK_posedge,
		TestSignal     => RADDR_ipd(4),
		TestSignalName => "RADDR(4)",
		TestDelay      => 0 ns,
		RefSignal      => RCLK_ipd,
		RefSignalName  => "RCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(4),
		SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(4),
		HoldLow        => thold_RADDR_RCLK_posedge_posedge(4),
		HoldHigh       => thold_RADDR_RCLK_negedge_posedge(4),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_RADDR5_RCLK_posedge,
		TimingData     => Tmkr_RADDR5_RCLK_posedge,
		TestSignal     => RADDR_ipd(5),
		TestSignalName => "RADDR(5)",
		TestDelay      => 0 ns,
		RefSignal      => RCLK_ipd,
		RefSignalName  => "RCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(5),
		SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(5),
		HoldLow        => thold_RADDR_RCLK_posedge_posedge(5),
		HoldHigh       => thold_RADDR_RCLK_negedge_posedge(5),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_RADDR6_RCLK_posedge,
		TimingData     => Tmkr_RADDR6_RCLK_posedge,
		TestSignal     => RADDR_ipd(6),
		TestSignalName => "RADDR(6)",
		TestDelay      => 0 ns,
		RefSignal      => RCLK_ipd,
		RefSignalName  => "RCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(6),
		SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(6),
		HoldLow        => thold_RADDR_RCLK_posedge_posedge(6),
		HoldHigh       => thold_RADDR_RCLK_negedge_posedge(6),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);


	      VitalSetupHoldCheck (
		Violation      => Tviol_RADDR7_RCLK_posedge,
		TimingData     => Tmkr_RADDR7_RCLK_posedge,
		TestSignal     => RADDR_ipd(7),
		TestSignalName => "RADDR(7)",
		TestDelay      => 0 ns,
		RefSignal      => RCLK_ipd,
		RefSignalName  => "RCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(7),
		SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(7),
		HoldLow        => thold_RADDR_RCLK_posedge_posedge(7),
		HoldHigh       => thold_RADDR_RCLK_negedge_posedge(7),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_RADDR8_RCLK_posedge,
		TimingData     => Tmkr_RADDR8_RCLK_posedge,
		TestSignal     => RADDR_ipd(8),
		TestSignalName => "RADDR(8)",
		TestDelay      => 0 ns,
		RefSignal      => RCLK_ipd,
		RefSignalName  => "RCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(8),
		SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(8),
		HoldLow        => thold_RADDR_RCLK_posedge_posedge(8),
		HoldHigh       => thold_RADDR_RCLK_negedge_posedge(8),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_RADDR9_RCLK_posedge,
		TimingData     => Tmkr_RADDR9_RCLK_posedge,
		TestSignal     => RADDR_ipd(9),
		TestSignalName => "RADDR(9)",
		TestDelay      => 0 ns,
		RefSignal      => RCLK_ipd,
		RefSignalName  => "RCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(9),
		SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(9),
		HoldLow        => thold_RADDR_RCLK_posedge_posedge(9),
		HoldHigh       => thold_RADDR_RCLK_negedge_posedge(9),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_RADDR10_RCLK_posedge,
		TimingData     => Tmkr_RADDR10_RCLK_posedge,
		TestSignal     => RADDR_ipd(10),
		TestSignalName => "RADDR(10)",
		TestDelay      => 0 ns,
		RefSignal      => RCLK_ipd,
		RefSignalName  => "RCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(10),
		SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(10),
		HoldLow        => thold_RADDR_RCLK_posedge_posedge(10),
		HoldHigh       => thold_RADDR_RCLK_negedge_posedge(10),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_RCLKE_RCLK_posedge,
		TimingData     => Tmkr_RCLKE_RCLK_posedge,
		TestSignal     => RCLKE_ipd,
		TestSignalName => "RCLKE",
		TestDelay      => 0 ns,
		RefSignal      => RCLK_ipd,
		RefSignalName  => "RCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_RCLKE_RCLK_posedge_posedge,
		SetupLow       => tsetup_RCLKE_RCLK_negedge_posedge,
		HoldLow        => thold_RCLKE_RCLK_posedge_posedge,
		HoldHigh       => thold_RCLKE_RCLK_negedge_posedge,
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_RE_RCLK_posedge,
		TimingData     => Tmkr_RE_RCLK_posedge,
		TestSignal     => RCLK_ipd,
		TestSignalName => "RCLK",
		TestDelay      => 0 ns,
		RefSignal      => RCLK_ipd,
		RefSignalName  => "RCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_RE_RCLK_posedge_posedge,
		SetupLow       => tsetup_RE_RCLK_negedge_posedge,
		HoldLow        => thold_RE_RCLK_posedge_posedge,
		HoldHigh       => thold_RE_RCLK_negedge_posedge,
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		       

	      VitalPeriodPulseCheck (
		Violation      => Pviol_RCLK,
		PeriodData     => PInfo_RCLK,
		TestSignal     => RCLK_ipd,
		TestSignalName => "RCLK",
		TestDelay      => 0 ns,
		Period         => 0 ns,
		PulseWidthHigh => tpw_RCLK_posedge,
		PulseWidthLow  => tpw_RCLK_negedge,
		CheckEnabled   => true,
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_WADDR0_WCLK_posedge,
		TimingData     => Tmkr_WADDR0_WCLK_posedge,
		TestSignal     => WADDR_ipd(0),
		TestSignalName => "WADDR(0)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(0),
		SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(0),
		HoldLow        => thold_WADDR_WCLK_posedge_posedge(0),
		HoldHigh       => thold_WADDR_WCLK_negedge_posedge(0),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_WADDR1_WCLK_posedge,
		TimingData     => Tmkr_WADDR1_WCLK_posedge,
		TestSignal     => WADDR_ipd(1),
		TestSignalName => "WADDR(1)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(1),
		SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(1),
		HoldLow        => thold_WADDR_WCLK_posedge_posedge(1),
		HoldHigh       => thold_WADDR_WCLK_negedge_posedge(1),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_WADDR2_WCLK_posedge,
		TimingData     => Tmkr_WADDR2_WCLK_posedge,
		TestSignal     => WADDR_ipd(2),
		TestSignalName => "WADDR(2)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(2),
		SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(2),
		HoldLow        => thold_WADDR_WCLK_posedge_posedge(2),
		HoldHigh       => thold_WADDR_WCLK_negedge_posedge(2),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_WADDR3_WCLK_posedge,
		TimingData     => Tmkr_WADDR3_WCLK_posedge,
		TestSignal     => WADDR_ipd(3),
		TestSignalName => "WADDR(3)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(3),
		SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(3),
		HoldLow        => thold_WADDR_WCLK_posedge_posedge(3),
		HoldHigh       => thold_WADDR_WCLK_negedge_posedge(3),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_WADDR4_WCLK_posedge,
		TimingData     => Tmkr_WADDR4_WCLK_posedge,
		TestSignal     => WADDR_ipd(4),
		TestSignalName => "WADDR(4)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(4),
		SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(4),
		HoldLow        => thold_WADDR_WCLK_posedge_posedge(4),
		HoldHigh       => thold_WADDR_WCLK_negedge_posedge(4),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_WADDR5_WCLK_posedge,
		TimingData     => Tmkr_WADDR5_WCLK_posedge,
		TestSignal     => WADDR_ipd(5),
		TestSignalName => "WADDR(5)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(5),
		SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(5),
		HoldLow        => thold_WADDR_WCLK_posedge_posedge(5),
		HoldHigh       => thold_WADDR_WCLK_negedge_posedge(5),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_WADDR6_WCLK_posedge,
		TimingData     => Tmkr_WADDR6_WCLK_posedge,
		TestSignal     => WADDR_ipd(6),
		TestSignalName => "WADDR(6)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(6),
		SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(6),
		HoldLow        => thold_WADDR_WCLK_posedge_posedge(6),
		HoldHigh       => thold_WADDR_WCLK_negedge_posedge(6),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_WADDR7_WCLK_posedge,
		TimingData     => Tmkr_WADDR7_WCLK_posedge,
		TestSignal     => WADDR_ipd(7),
		TestSignalName => "WADDR(7)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(7),
		SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(7),
		HoldLow        => thold_WADDR_WCLK_posedge_posedge(7),
		HoldHigh       => thold_WADDR_WCLK_negedge_posedge(7),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);


	      VitalSetupHoldCheck (
		Violation      => Tviol_WADDR8_WCLK_posedge,
		TimingData     => Tmkr_WADDR8_WCLK_posedge,
		TestSignal     => WADDR_ipd(8),
		TestSignalName => "WADDR(8)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(8),
		SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(8),
		HoldLow        => thold_WADDR_WCLK_posedge_posedge(8),
		HoldHigh       => thold_WADDR_WCLK_negedge_posedge(8),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);


	      VitalSetupHoldCheck (
		Violation      => Tviol_WADDR9_WCLK_posedge,
		TimingData     => Tmkr_WADDR9_WCLK_posedge,
		TestSignal     => WADDR_ipd(9),
		TestSignalName => "WADDR(9)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(9),
		SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(9),
		HoldLow        => thold_WADDR_WCLK_posedge_posedge(9),
		HoldHigh       => thold_WADDR_WCLK_negedge_posedge(9),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);


	      VitalSetupHoldCheck (
		Violation      => Tviol_WADDR10_WCLK_posedge,
		TimingData     => Tmkr_WADDR10_WCLK_posedge,
		TestSignal     => WADDR_ipd(10),
		TestSignalName => "WADDR(10)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(10),
		SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(10),
		HoldLow        => thold_WADDR_WCLK_posedge_posedge(10),
		HoldHigh       => thold_WADDR_WCLK_negedge_posedge(10),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_WCLKE_WCLK_posedge,
		TimingData     => Tmkr_WCLKE_WCLK_posedge,
		TestSignal     => WCLKE_ipd,
		TestSignalName => "WCLKE",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WCLKE_WCLK_posedge_posedge,
		SetupLow       => tsetup_WCLKE_WCLK_negedge_posedge,
		HoldLow        => thold_WCLKE_WCLK_posedge_posedge,
		HoldHigh       => thold_WCLKE_WCLK_negedge_posedge,
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_WE_WCLK_posedge,
		TimingData     => Tmkr_WE_WCLK_posedge,
		TestSignal     => WCLK_ipd,
		TestSignalName => "WCLK",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WE_WCLK_posedge_posedge,
		SetupLow       => tsetup_WE_WCLK_negedge_posedge,
		HoldLow        => thold_WE_WCLK_posedge_posedge,
		HoldHigh       => thold_WE_WCLK_negedge_posedge,
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	       VitalSetupHoldCheck (
		Violation      => Tviol_WDATA0_WCLK_posedge,
		TimingData     => Tmkr_WDATA0_WCLK_posedge,
		TestSignal     => WDATA_ipd(0),
		TestSignalName => "WDATA(0)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(0),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(0),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(0),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(0),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_WDATA1_WCLK_posedge,
		TimingData     => Tmkr_WDATA1_WCLK_posedge,
		TestSignal     => WDATA_ipd(1),
		TestSignalName => "WDATA(1)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(1),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(1),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(1),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(1),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_WDATA2_WCLK_posedge,
		TimingData     => Tmkr_WDATA2_WCLK_posedge,
		TestSignal     => WDATA_ipd(2),
		TestSignalName => "WDATA(2)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(2),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(2),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(2),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(2),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_WDATA3_WCLK_posedge,
		TimingData     => Tmkr_WDATA3_WCLK_posedge,
		TestSignal     => WDATA_ipd(3),
		TestSignalName => "WDATA(3)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(3),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(3),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(3),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(3),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_WDATA4_WCLK_posedge,
		TimingData     => Tmkr_WDATA4_WCLK_posedge,
		TestSignal     => WDATA_ipd(4),
		TestSignalName => "WDATA(4)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(4),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(4),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(4),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(4),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_WDATA5_WCLK_posedge,
		TimingData     => Tmkr_WDATA5_WCLK_posedge,
		TestSignal     => WDATA_ipd(5),
		TestSignalName => "WDATA(5)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(5),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(5),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(5),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(5),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_WDATA6_WCLK_posedge,
		TimingData     => Tmkr_WDATA6_WCLK_posedge,
		TestSignal     => WDATA_ipd(6),
		TestSignalName => "WDATA(6)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(6),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(6),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(6),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(6),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_WDATA7_WCLK_posedge,
		TimingData     => Tmkr_WDATA7_WCLK_posedge,
		TestSignal     => WDATA_ipd(7),
		TestSignalName => "WDATA(7)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(7),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(7),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(7),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(7),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	       VitalSetupHoldCheck (
		Violation      => Tviol_WDATA8_WCLK_posedge,
		TimingData     => Tmkr_WDATA8_WCLK_posedge,
		TestSignal     => WDATA_ipd(8),
		TestSignalName => "WDATA(8)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(8),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(8),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(8),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(8),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_WDATA9_WCLK_posedge,
		TimingData     => Tmkr_WDATA9_WCLK_posedge,
		TestSignal     => WDATA_ipd(9),
		TestSignalName => "WDATA(9)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(9),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(9),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(9),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(9),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_WDATA10_WCLK_posedge,
		TimingData     => Tmkr_WDATA10_WCLK_posedge,
		TestSignal     => WDATA_ipd(10),
		TestSignalName => "WDATA(10)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(10),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(10),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(10),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(10),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_WDATA11_WCLK_posedge,
		TimingData     => Tmkr_WDATA11_WCLK_posedge,
		TestSignal     => WDATA_ipd(11),
		TestSignalName => "WDATA(11)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(11),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(11),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(11),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(11),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_WDATA12_WCLK_posedge,
		TimingData     => Tmkr_WDATA12_WCLK_posedge,
		TestSignal     => WDATA_ipd(12),
		TestSignalName => "WDATA(12)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(12),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(12),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(12),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(12),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_WDATA13_WCLK_posedge,
		TimingData     => Tmkr_WDATA13_WCLK_posedge,
		TestSignal     => WDATA_ipd(13),
		TestSignalName => "WDATA(13)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(13),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(13),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(13),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(13),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_WDATA14_WCLK_posedge,
		TimingData     => Tmkr_WDATA14_WCLK_posedge,
		TestSignal     => WDATA_ipd(14),
		TestSignalName => "WDATA(14)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(14),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(14),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(14),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(14),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_WDATA15_WCLK_posedge,
		TimingData     => Tmkr_WDATA15_WCLK_posedge,
		TestSignal     => WDATA_ipd(15),
		TestSignalName => "WDATA(15)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(15),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(15),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(15),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(15),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	       VitalSetupHoldCheck (
		Violation      => Tviol_MASK0_WCLK_posedge,
		TimingData     => Tmkr_MASK0_WCLK_posedge,
		TestSignal     => MASK_ipd(0),
		TestSignalName => "MASK(0)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(0),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(0),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(0),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(0),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_MASK1_WCLK_posedge,
		TimingData     => Tmkr_MASK1_WCLK_posedge,
		TestSignal     => MASK_ipd(1),
		TestSignalName => "MASK(1)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(1),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(1),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(1),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(1),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_MASK2_WCLK_posedge,
		TimingData     => Tmkr_MASK2_WCLK_posedge,
		TestSignal     => MASK_ipd(2),
		TestSignalName => "MASK(2)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(2),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(2),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(2),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(2),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_MASK3_WCLK_posedge,
		TimingData     => Tmkr_MASK3_WCLK_posedge,
		TestSignal     => MASK_ipd(3),
		TestSignalName => "MASK(3)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(3),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(3),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(3),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(3),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_MASK4_WCLK_posedge,
		TimingData     => Tmkr_MASK4_WCLK_posedge,
		TestSignal     => MASK_ipd(4),
		TestSignalName => "MASK(4)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(4),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(4),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(4),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(4),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_MASK5_WCLK_posedge,
		TimingData     => Tmkr_MASK5_WCLK_posedge,
		TestSignal     => MASK_ipd(5),
		TestSignalName => "MASK(5)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(5),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(5),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(5),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(5),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_MASK6_WCLK_posedge,
		TimingData     => Tmkr_MASK6_WCLK_posedge,
		TestSignal     => MASK_ipd(6),
		TestSignalName => "MASK(6)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(6),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(6),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(6),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(6),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_MASK7_WCLK_posedge,
		TimingData     => Tmkr_MASK7_WCLK_posedge,
		TestSignal     => MASK_ipd(7),
		TestSignalName => "MASK(7)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(7),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(7),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(7),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(7),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	       VitalSetupHoldCheck (
		Violation      => Tviol_MASK8_WCLK_posedge,
		TimingData     => Tmkr_MASK8_WCLK_posedge,
		TestSignal     => MASK_ipd(8),
		TestSignalName => "MASK(8)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(8),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(8),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(8),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(8),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_MASK9_WCLK_posedge,
		TimingData     => Tmkr_MASK9_WCLK_posedge,
		TestSignal     => MASK_ipd(9),
		TestSignalName => "MASK(9)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(9),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(9),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(9),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(9),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_MASK10_WCLK_posedge,
		TimingData     => Tmkr_MASK10_WCLK_posedge,
		TestSignal     => MASK_ipd(10),
		TestSignalName => "MASK(10)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(10),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(10),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(10),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(10),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_MASK11_WCLK_posedge,
		TimingData     => Tmkr_MASK11_WCLK_posedge,
		TestSignal     => MASK_ipd(11),
		TestSignalName => "MASK(11)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(11),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(11),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(11),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(11),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_MASK12_WCLK_posedge,
		TimingData     => Tmkr_MASK12_WCLK_posedge,
		TestSignal     => MASK_ipd(12),
		TestSignalName => "MASK(12)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(12),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(12),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(12),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(12),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_MASK13_WCLK_posedge,
		TimingData     => Tmkr_MASK13_WCLK_posedge,
		TestSignal     => MASK_ipd(13),
		TestSignalName => "MASK(13)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(13),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(13),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(13),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(13),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_MASK14_WCLK_posedge,
		TimingData     => Tmkr_MASK14_WCLK_posedge,
		TestSignal     => MASK_ipd(14),
		TestSignalName => "MASK(14)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(14),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(14),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(14),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(14),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_MASK15_WCLK_posedge,
		TimingData     => Tmkr_MASK15_WCLK_posedge,
		TestSignal     => MASK_ipd(15),
		TestSignalName => "MASK(15)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(15),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(15),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(15),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(15),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
	   

	      VitalPeriodPulseCheck (
		Violation      => Pviol_WCLK,
		PeriodData     => PInfo_WCLK,
		TestSignal     => WCLK_ipd,
		TestSignalName => "WCLK",
		TestDelay      => 0 ns,
		Period         => 0 ns,
		PulseWidthHigh => tpw_WCLK_posedge,
		PulseWidthLow  => tpw_WCLK_negedge,
		CheckEnabled   => true,
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	    Violation  := Pviol_RCLK or
			  Tviol_RADDR0_RCLK_posedge or
			  Tviol_RADDR1_RCLK_posedge or
			  Tviol_RADDR2_RCLK_posedge or
			  Tviol_RADDR3_RCLK_posedge or
			  Tviol_RADDR4_RCLK_posedge or
			  Tviol_RADDR5_RCLK_posedge or
			  Tviol_RADDR6_RCLK_posedge or
			  Tviol_RADDR7_RCLK_posedge or
			  Tviol_RADDR8_RCLK_posedge or
			  Tviol_RADDR9_RCLK_posedge or
			  Tviol_RADDR10_RCLK_posedge or
			  Tviol_RCLKE_RCLK_posedge or
			  Tviol_RE_RCLK_posedge or
    			  Pviol_WCLK or
			  Tviol_WADDR0_WCLK_posedge or
			  Tviol_WADDR1_WCLK_posedge or
			  Tviol_WADDR2_WCLK_posedge or
			  Tviol_WADDR3_WCLK_posedge or
			  Tviol_WADDR4_WCLK_posedge or
			  Tviol_WADDR5_WCLK_posedge or
			  Tviol_WADDR6_WCLK_posedge or
			  Tviol_WADDR7_WCLK_posedge or
			  Tviol_WADDR8_WCLK_posedge or
			  Tviol_WADDR9_WCLK_posedge or
			  Tviol_WADDR10_WCLK_posedge or
			  Tviol_WCLKE_WCLK_posedge or
			  Tviol_WE_WCLK_posedge or
			  Tviol_WDATA0_WCLK_posedge or
			  Tviol_WDATA1_WCLK_posedge or
			  Tviol_WDATA2_WCLK_posedge or
			  Tviol_WDATA3_WCLK_posedge or
			  Tviol_WDATA4_WCLK_posedge or
			  Tviol_WDATA5_WCLK_posedge or
			  Tviol_WDATA6_WCLK_posedge or
			  Tviol_WDATA7_WCLK_posedge or
			  Tviol_WDATA8_WCLK_posedge or
			  Tviol_WDATA9_WCLK_posedge or
			  Tviol_WDATA10_WCLK_posedge or
			  Tviol_WDATA11_WCLK_posedge or
			  Tviol_WDATA12_WCLK_posedge or
			  Tviol_WDATA13_WCLK_posedge or
			  Tviol_WDATA14_WCLK_posedge or
			  Tviol_WDATA15_WCLK_posedge or
			  Tviol_MASK0_WCLK_posedge or
			  Tviol_MASK1_WCLK_posedge or
			  Tviol_MASK2_WCLK_posedge or
			  Tviol_MASK3_WCLK_posedge or
			  Tviol_MASK4_WCLK_posedge or
			  Tviol_MASK5_WCLK_posedge or
			  Tviol_MASK6_WCLK_posedge or
			  Tviol_MASK7_WCLK_posedge or
			  Tviol_MASK8_WCLK_posedge or
			  Tviol_MASK9_WCLK_posedge or
			  Tviol_MASK10_WCLK_posedge or
			  Tviol_MASK11_WCLK_posedge or
			  Tviol_MASK12_WCLK_posedge or
			  Tviol_MASK13_WCLK_posedge or
			  Tviol_MASK14_WCLK_posedge or
			  Tviol_MASK15_WCLK_posedge;

		assert violation = '0'
			report " Incorrect due to Timing Violations\n"
		severity warning;

	    end if ;
    end process TimingChecks;

------------------------
--  BEHAVIOR SECTION
------------------------

	READ_ADDR_HB <= RADDR_ipd(10) & RADDR_ipd(9) & RADDR_ipd(8);
	WRITE_ADDR_HB <= WADDR_ipd(10) & WADDR_ipd(9) & WADDR_ipd(8);
	READ_ADDR_LB <= RADDR_ipd(7) & RADDR_ipd(6) & RADDR_ipd(5)& RADDR_ipd(4) & RADDR_ipd(3) & RADDR_ipd(2) & RADDR_ipd(1) & RADDR_ipd(0);
	WRITE_ADDR_LB <= WADDR_ipd(7) & WADDR_ipd(6) & WADDR_ipd(5)& WADDR_ipd(4) & WADDR_ipd(3) & WADDR_ipd(2) & WADDR_ipd(1) & WADDR_ipd(0);

	LatchAddress:process(RCLK_ipd) 
	begin 
		if(RCLK_ipd'event and RCLK_ipd='1') then 
		READ_ADDR_HB_reg <=READ_ADDR_HB;  
		end if; 
	end process LatchAddress;   

	read_data_decoder_inst  : read_data_decoder 
		generic map (
			READ_MODE => READ_MODE
		)
		port map (
			di	=> RD,
			ai	=> READ_ADDR_HB_reg,
			ldo	=> RDATA_zd
		);

	
	write_data_decoder_inst  : write_data_decoder
		generic map (
			WRITE_MODE => WRITE_MODE
		)
		port map (
			di  => WDATA_ipd,
			ldo  => WD
		);

	mask_data_decoder_inst : mask_decoder
		generic map (
			WRITE_MODE => WRITE_MODE
		)
		port map (
			mi  => MASK_ipd,
			mo  => MASK_RAM,
			ai  => WRITE_ADDR_HB
		);
	ram_inst : SB_RAM4K
		generic map (
			INIT_0     => INIT_0,
			INIT_1     => INIT_1,
			INIT_2     => INIT_2,
			INIT_3     => INIT_3,
			INIT_4     => INIT_4,
			INIT_5     => INIT_5,
			INIT_6     => INIT_6,
			INIT_7     => INIT_7,
			INIT_8     => INIT_8,
			INIT_9     => INIT_9,
			INIT_A     => INIT_A,
			INIT_B     => INIT_B,
			INIT_C     => INIT_C,
			INIT_D     => INIT_D,
			INIT_E     => INIT_E,
			INIT_F     => INIT_F
		)
		port map (
			RDATA	=> RD,
			RCLK	=> RCLK_ipd,
			RCLKE	=> RCLKE_ipd,
			RE	=> RE_ipd,
			RADDR	=> READ_ADDR_LB,
			MASK	=> MASK_RAM,
			WDATA	=> WD,       
			WCLK	=> WCLK_ipd,
			WCLKE	=> WCLKE_ipd,
			WE	=> WE_ipd,
			WADDR	=> WRITE_ADDR_LB
		);

------------------------
--  Path Delay Section
------------------------
	PathDelay : process(RDATA_zd)

	variable RDATA_GlitchData0  : VitalGlitchDataType;
	variable RDATA_GlitchData1  : VitalGlitchDataType;
	variable RDATA_GlitchData2  : VitalGlitchDataType;
	variable RDATA_GlitchData3  : VitalGlitchDataType;
	variable RDATA_GlitchData4  : VitalGlitchDataType;
	variable RDATA_GlitchData5  : VitalGlitchDataType;
	variable RDATA_GlitchData6  : VitalGlitchDataType;
	variable RDATA_GlitchData7  : VitalGlitchDataType;
	variable RDATA_GlitchData8  : VitalGlitchDataType;
	variable RDATA_GlitchData9  : VitalGlitchDataType;
	variable RDATA_GlitchData10 : VitalGlitchDataType;
	variable RDATA_GlitchData11 : VitalGlitchDataType;
	variable RDATA_GlitchData12 : VitalGlitchDataType;
	variable RDATA_GlitchData13 : VitalGlitchDataType;
	variable RDATA_GlitchData14 : VitalGlitchDataType;
	variable RDATA_GlitchData15 : VitalGlitchDataType;
	begin
	    VitalPathDelay01 (
	      OutSignal     => RDATA(0),
	      GlitchData    => RDATA_GlitchData0,
	      OutSignalName => "RDATA(0)",
	      OutTemp       => RDATA_zd(0),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(0), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => RDATA(1),
	      GlitchData    => RDATA_GlitchData1,
	      OutSignalName => "RDATA(1)",
	      OutTemp       => RDATA_zd(1),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(1), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => RDATA(2),
	      GlitchData    => RDATA_GlitchData2,
	      OutSignalName => "RDATA(2)",
	      OutTemp       => RDATA_zd(2),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(2), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => RDATA(3),
	      GlitchData    => RDATA_GlitchData3,
	      OutSignalName => "RDATA(3)",
	      OutTemp       => RDATA_zd(3),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(3), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => RDATA(4),
	      GlitchData    => RDATA_GlitchData4,
	      OutSignalName => "RDATA(4)",
	      OutTemp       => RDATA_zd(4),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(4), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => RDATA(5),
	      GlitchData    => RDATA_GlitchData5,
	      OutSignalName => "RDATA(5)",
	      OutTemp       => RDATA_zd(5),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(5), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => RDATA(6),
	      GlitchData    => RDATA_GlitchData6,
	      OutSignalName => "RDATA(6)",
	      OutTemp       => RDATA_zd(6),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(6), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => RDATA(7),
	      GlitchData    => RDATA_GlitchData7,
	      OutSignalName => "RDATA(7)",
	      OutTemp       => RDATA_zd(7),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(7), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => RDATA(8),
	      GlitchData    => RDATA_GlitchData8,
	      OutSignalName => "RDATA(8)",
	      OutTemp       => RDATA_zd(8),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(8), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => RDATA(9),
	      GlitchData    => RDATA_GlitchData9,
	      OutSignalName => "RDATA(9)",
	      OutTemp       => RDATA_zd(9),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(9), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => RDATA(10),
	      GlitchData    => RDATA_GlitchData10,
	      OutSignalName => "RDATA(10)",
	      OutTemp       => RDATA_zd(10),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(10), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => RDATA(11),
	      GlitchData    => RDATA_GlitchData11,
	      OutSignalName => "RDATA(11)",
	      OutTemp       => RDATA_zd(11),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(11), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => RDATA(12),
	      GlitchData    => RDATA_GlitchData12,
	      OutSignalName => "RDATA(12)",
	      OutTemp       => RDATA_zd(12),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(12), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => RDATA(13),
	      GlitchData    => RDATA_GlitchData13,
	      OutSignalName => "RDATA(13)",
	      OutTemp       => RDATA_zd(13),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(13), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => RDATA(14),
	      GlitchData    => RDATA_GlitchData14,
	      OutSignalName => "RDATA(14)",
	      OutTemp       => RDATA_zd(14),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(14), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => RDATA(15),
	      GlitchData    => RDATA_GlitchData15,
	      OutSignalName => "RDATA(15)",
	      OutTemp       => RDATA_zd(15),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(15), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	end process;

	end block;


end SB_RAM40_4K_V;   --- SB_RAM40_4K


library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity read_data_decoder is
	generic (
		READ_MODE : integer := 0
	);
	port (
	 	di  : in std_logic_vector (15 downto 0);
		ldo  : out std_logic_vector (15 downto 0);
		ai  : in std_logic_vector (2 downto 0)
	);
end read_data_decoder;

architecture read_data_decoder_arch of read_data_decoder is
	signal mode : std_logic_vector ( 1 downto 0);
	signal selector : std_logic_vector (4 downto 0);
begin
	selector <= mode & ai;

	process
	begin
		if(READ_MODE = 0)
		then
			mode <= "00";
		else
			if(READ_MODE = 1)
			then
				mode <= "01";
			else
				if(READ_MODE = 2)
				then
					mode <= "10";
				else
					if(READ_MODE = 3)
					then
						mode <=  "11";
					else
						assert false
						report "SBT ERROR: Unknown RAM modes\n Valid modes are 0 (256X16), 1 (512X8), 2 (1024X4), 3 (2048X2)\n"
						severity error;
					end if;
				end if;
			end if;
		end if;
		wait;
	end process;

	process (selector, di ) 
	begin
		case selector is
			when "00000" | "00001" | "00010" | "00011" | "00100"| "00101" | "00110" | "00111" => 
				ldo <= di;
			when "01000" | "01010" | "01100" | "01110" => 
				ldo <= '0' & di(14) & '0' & di(12) &'0' & di(10) &'0' & di(8) &'0' & di(6) &'0' & di(4) &'0' & di(2) &'0' & di(0) ;
			when "01001" | "01011" | "01101" | "01111" => 
				ldo <= '0' & di(15) & '0' & di(13) &'0' & di(11) &'0' & di(9) &'0' & di(7) &'0' & di(5) &'0' & di(3) &'0' & di(1) ;
			when "10000" | "10100" =>
				ldo <= "00" & di(12) & "000" & di(8) & "000" &  di(4) & "000" & di(0) & "0" ;
			when "10001" | "10101" =>
				ldo <= "00" & di(13) & "000" & di(9) & "000" &  di(5) & "000" & di(1) & "0" ;
			when "10010" | "10110" =>
				ldo <= "00" & di(14) & "000" & di(10) & "000" &  di(6) & "000" & di(2) & "0" ;
			when "10011" | "10111" =>
				ldo <= "00" & di(15) & "000" & di(11) & "000" &  di(7) & "000" & di(3) & "0" ;
			when "11000" =>
				ldo <= "0000" & di(8) & "0000000" & di(0) & "000";
			when "11001" =>
				ldo <= "0000" & di(9) & "0000000" & di(1) & "000";
			when "11010" =>
				ldo <= "0000" & di(10) & "0000000" & di(2) & "000";
			when "11011" =>
				ldo <= "0000" & di(11) & "0000000" & di(3) & "000";
			when "11100" =>
				ldo <= "0000" & di(12) & "0000000" & di(4) & "000";
			when "11101" =>
				ldo <= "0000" & di(13) & "0000000" & di(5) & "000";
			when "11110" =>
				ldo <= "0000" & di(14) & "0000000" & di(6) & "000";
			when "11111" =>
				ldo <= "0000" & di(15) & "0000000" & di(7) & "000";
			when others => 
			--	assert false
			        assert (NOW=0 ns) or (NOW = 0 ps) 	
				report "SBT ERROR: End up in unknown State during Read data decoding. If this occurs at zero simulation time (0ps/0ns) this error msg can be ignored \n"
				severity error;
		end case;
	end process;
end read_data_decoder_arch;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity write_data_decoder is
	generic (
		WRITE_MODE : integer := 0
	);
	port (
	 	di  : in std_logic_vector (15 downto 0);
		ldo  : out std_logic_vector (15 downto 0)
	);
end write_data_decoder;

architecture write_data_decoder_arch of write_data_decoder is
	signal mode : std_logic_vector ( 1 downto 0);
	signal selector : std_logic_vector (1 downto 0);
begin
	selector <= mode ;

	process
	begin
		if(WRITE_MODE = 0)
		then
			mode <= "00";
		else
			if(WRITE_MODE = 1)
			then
				mode <= "01";
			else
				if(WRITE_MODE = 2)
				then
					mode <= "10";
				else
					if(WRITE_MODE = 3)
					then
						mode <=  "11";
					else
						assert false
						report "SBT ERROR: Unknown RAM modes\n Valid modes are 0 (256X16), 1 (512X8), 2 (1024X4), 3 (2048X2)\n"
						severity error;
					end if;
				end if;
			end if;
		end if;
		wait;
	end process;

	process (selector, di )
	begin
		case selector is
			when "00" => 
				ldo <= di;
			when "01" => 
				ldo <= di(14) & di(14) & di(12) & di(12) & di(10) & di(10) & di(8) & di(8) & di(6) & di(6) & di(4) & di(4) & di(2) & di(2) & di(0) & di(0) ; 
			when "10" => 
				ldo <= di(13) & di(13) & di(13) & di(13) & di(9) & di(9) & di(9) & di(9) & di(5) & di(5) & di(5) & di(5) & di(1) & di(1) & di(1) & di(1) ; 
			when "11" =>
				ldo <= di(11) & di(11) & di(11) & di(11) & di(11) & di(11) & di(11) & di(11) & di(3) & di(3) & di(3) & di(3) & di(3) & di(3) & di(3) & di(3) ; 
			when others => 
			--	assert false
				assert (NOW=0 ns) or (NOW = 0 ps)		
				report "SBT ERROR : End up in unknown State during write data decoding. If this occurs at zero simulation time (0ps/0ns) this can be ignored\n"
				severity error;
		end case;
	end process;
end write_data_decoder_arch;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity mask_decoder is
	generic (
		WRITE_MODE : integer := 0
	);
	port (
	 	mi  : in std_logic_vector (15 downto 0);
		mo  : out std_logic_vector (15 downto 0);
		ai  : in std_logic_vector (2 downto 0)
	);
end mask_decoder;

architecture mask_data_decoder_arch of mask_decoder is
	signal mode : std_logic_vector ( 1 downto 0);
	signal selector : std_logic_vector (4 downto 0);
begin
	selector <= mode & ai;

	process
	begin
		if(WRITE_MODE = 0)
		then
			mode <= "00";
		else
			if(WRITE_MODE = 1)
			then
				mode <= "01";
			else
				if(WRITE_MODE = 2)
				then
					mode <= "10";
				else
					if(WRITE_MODE = 3)
					then
						mode <=  "11";
					else
						assert false
						report "SBT ERROR: Unknown RAM modes\n Valid modes are 256X16, 512X8, 1024X4, 2048X2\n"
						severity error;
					end if;
				end if;
			end if;
		end if;
		wait;
	end process;

	process (selector, mi )
	begin
		case selector is
			when "00000" | "00001" | "00010" | "00011" | "00100"| "00101" | "00110" | "00111" => 
				mo <= mi;
			when "01000" | "01010" | "01100" | "01110" => 
				mo <= X"AAAA";
			when "01001" | "01011" | "01101" | "01111" => 
				mo <= X"5555";
			when "10000" | "10100" =>
				mo <= X"EEEE";
			when "10001" | "10101" =>
				mo <= X"DDDD";
			when "10010" | "10110" =>
				mo <= X"BBBB";
			when "10011" | "10111" =>
				mo <= X"7777";
			when "11000" =>
				mo <= X"FEFE";
			when "11001" =>
				mo <= X"FDFD";
			when "11010" =>
				mo <= X"FBFB";
			when "11011" =>
				mo <= X"F7F7";
			when "11100" =>
				mo <= X"EFEF";
			when "11101" =>
				mo <= X"DFDF";
			when "11110" =>
				mo <= X"BFBF";
			when "11111" =>
				mo <= X"7F7F";
			when others => 				
			--	assert false
				assert (NOW=0 ns) or (NOW = 0 ps)		
				report "SBT ERROR : End up in unknown State during mask data decoding. If this occurs at zero simulation time (0ps/0ns) this can be ignored \n"
				severity error;
		end case;
	end process;
end mask_data_decoder_arch;

---------------------------------------
	--- SB_RAM40_4KNR
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM40_4KNR is

  generic ( 
  	   WRITE_MODE : integer := 0; -- can be integer 0(256X16 mode) or 1(512X8 mode) or 2(1024X4 mode) or 3(2048X2 mode)
  	   READ_MODE  : integer := 0; -- can be integer 0(256X16 mode) or 1(512X8 mode) or 2(1024X4 mode) or 3(2048X2 mode)
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 15  downto 0) ;
                RCLKN : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'L';
                RADDR : in  std_logic_vector( 10  downto 0) ;
                WCLK  : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'L';
                WADDR : in  std_logic_vector( 10  downto 0) ;
                MASK  : in  std_logic_vector( 15  downto 0) ;
                WDATA : in  std_logic_vector( 15 downto 0)
               );
  
  
end SB_RAM40_4KNR;

architecture SB_RAM40_4KNR_V of SB_RAM40_4KNR is
	component SB_RAM40_4K
		generic (
			WRITE_MODE : integer;
			READ_MODE  : integer;
			INIT_0	   : bit_vector;
			INIT_1	   : bit_vector;
			INIT_2	   : bit_vector;
			INIT_3	   : bit_vector;
			INIT_4	   : bit_vector;
			INIT_5	   : bit_vector;
			INIT_6	   : bit_vector;
			INIT_7	   : bit_vector;
			INIT_8	   : bit_vector;
			INIT_9	   : bit_vector;
			INIT_A	   : bit_vector;
			INIT_B	   : bit_vector;
			INIT_C	   : bit_vector;
			INIT_D	   : bit_vector;
			INIT_E	   : bit_vector;
			INIT_F	   : bit_vector
		);
		port (
			RDATA	   : out std_logic_vector(15 downto 0);
			RCLK	   : in std_logic;
			RCLKE	   : in std_logic;
			RE	   : in std_logic;
			RADDR	   : in std_logic_vector(10 downto 0);
			MASK	   : in std_logic_vector(15 downto 0);
			WDATA	   : in std_logic_vector(15 downto 0);
			WCLK	   : in std_logic;
			WCLKE	   : in std_logic;
			WE	   : in std_logic;
			WADDR	   : in std_logic_vector(10 downto 0)
		);
	end component;

	signal RCLK : std_logic;

begin
	RCLK <= not(RCLKN);
	ram40_4k_nr_inst : SB_RAM40_4K
		generic map (
			WRITE_MODE => WRITE_MODE,
			READ_MODE  => READ_MODE,
			INIT_0     => INIT_0,
			INIT_1     => INIT_1,
			INIT_2     => INIT_2,
			INIT_3     => INIT_3,
			INIT_4     => INIT_4,
			INIT_5     => INIT_5,
			INIT_6     => INIT_6,
			INIT_7     => INIT_7,
			INIT_8     => INIT_8,
			INIT_9     => INIT_9,
			INIT_A     => INIT_A,
			INIT_B     => INIT_B,
			INIT_C     => INIT_C,
			INIT_D     => INIT_D,
			INIT_E     => INIT_E,
			INIT_F     => INIT_F
		)
		port map (
			RDATA	=> RDATA,
			RCLK	=> RCLK,
			RCLKE	=> RCLKE,
			RE	=> RE,
			RADDR	=> RADDR,
			MASK	=> MASK,
			WDATA	=> WDATA,
			WCLK	=> WCLK,
			WCLKE	=> WCLKE,
			WE	=> WE,
			WADDR	=> WADDR
		);
end SB_RAM40_4KNR_V;   --- SB_RAM40_4KNR


---------------------------------------
	--- SB_RAM40_4KNW
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM40_4KNW is

  generic ( 
  	   WRITE_MODE : integer := 0; -- can be integer 0(256X16 mode) or 1(512X8 mode) or 2(1024X4 mode) or 3(2048X2 mode)
  	   READ_MODE  : integer := 0; -- can be integer 0(256X16 mode) or 1(512X8 mode) or 2(1024X4 mode) or 3(2048X2 mode)
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 15  downto 0) ;
                RCLK  : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'L';
                RADDR : in  std_logic_vector( 10  downto 0) ;
                WCLKN : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'L';
                WADDR : in  std_logic_vector( 10  downto 0) ;
                MASK  : in  std_logic_vector( 15  downto 0) ;
                WDATA : in  std_logic_vector( 15 downto 0)
               );
  
  
end SB_RAM40_4KNW;

architecture SB_RAM40_4KNW_V of SB_RAM40_4KNW is
	component SB_RAM40_4K
		generic (
			WRITE_MODE : integer;
			READ_MODE  : integer;
			INIT_0	   : bit_vector;
			INIT_1	   : bit_vector;
			INIT_2	   : bit_vector;
			INIT_3	   : bit_vector;
			INIT_4	   : bit_vector;
			INIT_5	   : bit_vector;
			INIT_6	   : bit_vector;
			INIT_7	   : bit_vector;
			INIT_8	   : bit_vector;
			INIT_9	   : bit_vector;
			INIT_A	   : bit_vector;
			INIT_B	   : bit_vector;
			INIT_C	   : bit_vector;
			INIT_D	   : bit_vector;
			INIT_E	   : bit_vector;
			INIT_F	   : bit_vector
		);
		port (
			RDATA	   : out std_logic_vector(15 downto 0);
			RCLK	   : in std_logic;
			RCLKE	   : in std_logic;
			RE	   : in std_logic;
			RADDR	   : in std_logic_vector(10 downto 0);
			MASK	   : in std_logic_vector(15 downto 0);
			WDATA	   : in std_logic_vector(15 downto 0);
			WCLK	   : in std_logic;
			WCLKE	   : in std_logic;
			WE	   : in std_logic;
			WADDR	   : in std_logic_vector(10 downto 0)
		);
	end component;

	signal WCLK : std_logic;

begin
	WCLK <= not(WCLKN);
	ram40_4k_nr_inst : SB_RAM40_4K
		generic map (
			WRITE_MODE => WRITE_MODE,
			READ_MODE  => READ_MODE,
			INIT_0     => INIT_0,
			INIT_1     => INIT_1,
			INIT_2     => INIT_2,
			INIT_3     => INIT_3,
			INIT_4     => INIT_4,
			INIT_5     => INIT_5,
			INIT_6     => INIT_6,
			INIT_7     => INIT_7,
			INIT_8     => INIT_8,
			INIT_9     => INIT_9,
			INIT_A     => INIT_A,
			INIT_B     => INIT_B,
			INIT_C     => INIT_C,
			INIT_D     => INIT_D,
			INIT_E     => INIT_E,
			INIT_F     => INIT_F
		)
		port map (
			RDATA	=> RDATA,
			RCLK	=> RCLK,
			RCLKE	=> RCLKE,
			RE	=> RE,
			RADDR	=> RADDR,
			MASK	=> MASK,
			WDATA	=> WDATA,
			WCLK	=> WCLK,
			WCLKE	=> WCLKE,
			WE	=> WE,
			WADDR	=> WADDR
		);
end SB_RAM40_4KNW_V;   --- SB_RAM40_4KNW


---------------------------------------
	--- SB_RAM40_4KNRNW
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM40_4KNRNW is

  generic ( 
  	   WRITE_MODE : integer := 0 ; -- can be integer 0(256X16 mode) or 1(512X8 mode) or 2(1024X4 mode) or 3(2048X2 mode)
  	   READ_MODE  : integer := 0 ; -- can be integer 0(256X16 mode) or 1(512X8 mode) or 2(1024X4 mode) or 3(2048X2 mode)
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 15  downto 0) ;
                RCLKN : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'L';
                RADDR : in  std_logic_vector( 10  downto 0) ;
                WCLKN : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'L';
                WADDR : in  std_logic_vector( 10  downto 0) ;
                MASK  : in  std_logic_vector( 15  downto 0) ;
                WDATA : in  std_logic_vector( 15 downto 0)
               );
  
  
end SB_RAM40_4KNRNW;

architecture SB_RAM40_4KNRNW_V of SB_RAM40_4KNRNW is
	component SB_RAM40_4K
		generic (
			WRITE_MODE : integer;
			READ_MODE  : integer;
			INIT_0	   : bit_vector;
			INIT_1	   : bit_vector;
			INIT_2	   : bit_vector;
			INIT_3	   : bit_vector;
			INIT_4	   : bit_vector;
			INIT_5	   : bit_vector;
			INIT_6	   : bit_vector;
			INIT_7	   : bit_vector;
			INIT_8	   : bit_vector;
			INIT_9	   : bit_vector;
			INIT_A	   : bit_vector;
			INIT_B	   : bit_vector;
			INIT_C	   : bit_vector;
			INIT_D	   : bit_vector;
			INIT_E	   : bit_vector;
			INIT_F	   : bit_vector
		);
		port (
			RDATA	   : out std_logic_vector(15 downto 0);
			RCLK	   : in std_logic;
			RCLKE	   : in std_logic;
			RE	   : in std_logic;
			RADDR	   : in std_logic_vector(10 downto 0);
			MASK	   : in std_logic_vector(15 downto 0);
			WDATA	   : in std_logic_vector(15 downto 0);
			WCLK	   : in std_logic;
			WCLKE	   : in std_logic;
			WE	   : in std_logic;
			WADDR	   : in std_logic_vector(10 downto 0)
		);
	end component;

	signal RCLK : std_logic;
	signal WCLK : std_logic;

begin
	RCLK <= not(RCLKN);
	WCLK <= not(WCLKN);
	ram40_4k_nr_inst : SB_RAM40_4K
		generic map (
			WRITE_MODE => WRITE_MODE,
			READ_MODE  => READ_MODE,
			INIT_0     => INIT_0,
			INIT_1     => INIT_1,
			INIT_2     => INIT_2,
			INIT_3     => INIT_3,
			INIT_4     => INIT_4,
			INIT_5     => INIT_5,
			INIT_6     => INIT_6,
			INIT_7     => INIT_7,
			INIT_8     => INIT_8,
			INIT_9     => INIT_9,
			INIT_A     => INIT_A,
			INIT_B     => INIT_B,
			INIT_C     => INIT_C,
			INIT_D     => INIT_D,
			INIT_E     => INIT_E,
			INIT_F     => INIT_F
		)
		port map (
			RDATA	=> RDATA,
			RCLK	=> RCLK,
			RCLKE	=> RCLKE,
			RE	=> RE,
			RADDR	=> RADDR,
			MASK	=> MASK,
			WDATA	=> WDATA,
			WCLK	=> WCLK,
			WCLKE	=> WCLKE,
			WE	=> WE,
			WADDR	=> WADDR
		);
end SB_RAM40_4KNRNW_V;   --- SB_RAM40_4KNRNW

--///////////////////////////////////// ---
	---  END ICE40 RAM Primitives ---
--///////////////////////////////////// ---

--------------------------------------------------------------------------
----- 		mux4to1 					    ---- 
--------------------------------------------------------------------------
--
--library IEEE;
--use IEEE.std_logic_1164.all;
--use IEEE.std_logic_arith.all;
--use IEEE.std_logic_unsigned.all;
--use IEEE.VITAL_Primitives.all;
--use IEEE.VITAL_Timing.all;
--use work.std_logic_SBT.all;
-- 
--
--entity  mux4to1   is
--	port ( 
--		a,b,c,d : in std_logic; 
--		sel 	: in std_logic_vector(1 downto 0); 
--		o	: out std_logic 
--	      ); 
--end mux4to1;
--
--
--architecture mux4to1_arch of mux4to1 is 
--begin  
--	process( a,b,c,d,sel) 
--	begin 
--	case(sel) is 
--		when "00" => o<=a; 
--		when "01" => o<=b; 
--		when "10" => o<=c; 
--		when "11" => o<=d; 
--		when others => o<='0'; 
--	end case; 
--  	end process; 
--end mux4to1_arch; 


------------------------------------------------------------------------
--- 		Delay4Buf				    ---- 
------------------------------------------------------------------------
--
--library IEEE;
--use IEEE.std_logic_1164.all;
--use IEEE.std_logic_arith.all;
--use IEEE.std_logic_unsigned.all;
--use IEEE.VITAL_Primitives.all;
--use IEEE.VITAL_Timing.all;
--use work.std_logic_SBT.all;
-- 
--
--entity Delay4Buf  is
--	generic ( 
--		BUF_DELAY       : time := 150 ps ; 
-- 		MUXINV_DELAY    : time := 0 ps
--		); 	
--	port  ( 
--		a 		:in std_logic;   	
--	 	s		:in std_logic_vector(1 downto 0); 
--		delay4bufout	:out std_logic; 
--		muxinvout	:out std_logic
--	       );   		
--end Delay4Buf;
--
--architecture Delay4Buf_arch of Delay4Buf is 
--
--component  mux4to1   is
--	port ( 
--		a,b,c,d : in std_logic; 
--		sel 	: in std_logic_vector(1 downto 0); 
--		o	: out std_logic 
--	      ); 
--end component ;
--
--signal buf1out, buf2out,buf3out, buf4out  : std_logic; 
--signal muxout 				  : std_logic; 
--begin 
--	-- delay tap
--	buf1out  <= a after BUF_DELAY; 	 
--	buf2out  <= buf1out  after BUF_DELAY; 
--	buf3out  <= buf2out  after BUF_DELAY; 
--	buf4out  <= buf3out  after BUF_DELAY ; 
--	
--	delay4bufout <= buf4out; 	       
--	
--	mux4to1_inst : mux4to1 
--	port map (
--		 a=>buf1out,
--		 b=>buf2out,
--		 c=>buf3out,
--		 d=>buf4out,
--		 sel=>s,
--		 o=>muxout
--		);   
--
--
----	muxinvout  <= not(muxout) after MUXINV_DELAY;     -- check 
--	muxinvout  <= not(muxout); 
--	
--end Delay4Buf_arch;  


------------------------------------------------------------------------
--- 		FineDlyAdj 					    ---- 
------------------------------------------------------------------------

--library IEEE;
--use IEEE.std_logic_1164.all;
--use IEEE.std_logic_arith.all;
--use IEEE.std_logic_unsigned.all;
--use IEEE.VITAL_Primitives.all;
--use IEEE.VITAL_Timing.all;
--use work.std_logic_SBT.all;
-- 
--
--entity FineDlyAdj  is
--	generic (
--		FIXED_DELAY_ADJUSTMENT   : bit_vector(3 downto 0) :="0000"; 
--		DELAY_ADJUSTMENT_MODE    : string 		  :="FIXED";
--		BUF_DELAY		 : time 		  := 150 ps;
--		MUXINV_DELAY		 : time 		  := 0 ps ); 
--	port 	( 
--		signalin		:in  std_logic; 
--		DlyAdj			:in  std_logic_vector(3 downto 0); 
--		delayedout 		:out std_logic
--		); 
--
--end FineDlyAdj; 
--
--architecture FineDlyAdj_arch of FineDlyAdj is 
--
--component Delay4Buf  is
--	generic ( 
--		BUF_DELAY       : time := 150 ps ; 
-- 		MUXINV_DELAY    : time := 0 ps
--		); 	
--	port  ( 
--		a 		:in std_logic;   	
--	 	s		:in std_logic_vector(1 downto 0); 
--		delay4bufout	:out std_logic; 
--		muxinvout	:out std_logic
--	       );   		
--end component; 
--
--component  mux4to1   is
--	port ( 
--		a,b,c,d : in std_logic; 
--		sel 	: in std_logic_vector(1 downto 0); 
--		o	: out std_logic 
--	      ); 
--end component ;
--
-- signal fixed_delay_adj_generic : std_logic_vector( 3 downto 0);
-- signal bufcntselector   	: std_logic_vector( 3 downto 0);  
-- signal delay4bufout1,delay4bufout2, delay4bufout3, delay4bufout4 : std_logic; 
-- signal muxinvout1, muxinvout2,muxinvout3,muxinvout4 : std_logic;  
-- signal l2muxout		: std_logic;
-- 
--begin 
--
-- -- generics
--	fixed_delay_adj_generic <= TO_STDLOGICVECTOR(FIXED_DELAY_ADJUSTMENT); 
-- 
-- -- validations -- Process with wait statement 
-- initial_proc :   process 
-- begin 
--
--  if (DELAY_ADJUSTMENT_MODE = "FIXED" and  (FIXED_DELAY_ADJUSTMENT > "1111" or  FIXED_DELAY_ADJUSTMENT < "0000" )) then 
--            report  ("************************SBT: ERROR ****************************");
--            report  ("Valid values for FIXED_DELAY_ADJUSTMENT parameter are 4'b0000 through 4'b1111");
--            report  ("Due to incorrect configuration of the PLL, the simulation results are invalid.");
--  end if; 	
--  if ((DELAY_ADJUSTMENT_MODE = "DYNAMIC") and (FIXED_DELAY_ADJUSTMENT /= "0000")) then 
--            report ("************************SBT: Info*****************************");
--            report ("Since DELAY_ADJUSTMENT_MODE=DYNAMIC, parameter FIXED_DELAY_ADJUSTMENT will be ignored.");
--            report ("Set FIXED_DELAY_ADJUSTMENT=0 to disable this message.");
--  end if ; 	
-- wait; 	-- wait forever 		
-- end process initial_proc; 	
--
-- 
-- -- logics 
-- process (DlyAdj,fixed_delay_adj_generic) 
-- begin 
--	if(DELAY_ADJUSTMENT_MODE = "FIXED") then 
--		bufcntselector <= fixed_delay_adj_generic ; 
--	else 
--		bufcntselector <= DlyAdj; 
--	end if ; 
-- end process;  
--
--
-- delay4bufinst1  : Delay4Buf
-- generic map ( 
--	  BUF_DELAY => BUF_DELAY, 
--	  MUXINV_DELAY => MUXINV_DELAY		
--	  ) 	
-- port map ( 
--	 a => signalin, 
--	 s => bufcntselector(1 downto 0), 
--	 delay4bufout => delay4bufout1,	
--	 muxinvout    => muxinvout1	
--	  ); 
--   		
--  
-- delay4bufinst2  : Delay4Buf
-- generic map ( 
--	  BUF_DELAY => BUF_DELAY, 
--	  MUXINV_DELAY => MUXINV_DELAY		
--	  ) 	
-- port map ( 
--	 a => delay4bufout1,  
--	 s => bufcntselector(1 downto 0), 
--	 delay4bufout => delay4bufout2,	
--	 muxinvout    => muxinvout2	
--	  ); 
-- 
-- delay4bufinst3  : Delay4Buf
-- generic map ( 
--	  BUF_DELAY => BUF_DELAY, 
--	  MUXINV_DELAY => MUXINV_DELAY		
--	  ) 	
-- port map ( 
--	 a => delay4bufout2, 
--	 s => bufcntselector(1 downto 0), 
--	 delay4bufout => delay4bufout3,	
--	 muxinvout    => muxinvout3	
--	  ); 
--
-- delay4bufinst4  : Delay4Buf
-- generic map ( 
--	  BUF_DELAY => BUF_DELAY, 
--	  MUXINV_DELAY => MUXINV_DELAY		
--	  ) 	
-- port map ( 
--	 a => delay4bufout3,  
--	 s => bufcntselector(1 downto 0), 
--	 delay4bufout => delay4bufout4,	
--	 muxinvout    => muxinvout4	
--	  ); 
--
--
--  mux4to1_level2 : mux4to1 
--	port map (
--		 a=>muxinvout1,
--		 b=>muxinvout2,
--		 c=>muxinvout3,
--		 d=>muxinvout4,
--		 sel=>bufcntselector(3 downto 2),
--		 o=>l2muxout
--		);   
--
----	delayedout <= l2muxout after MUXINV_DELAY; 	
--	delayedout <= not(l2muxout) after MUXINV_DELAY; 
--	
--end FineDlyAdj_arch; 
--
--
--------------------------------------------------------
------ 		ShiftReg427 			  ---- 
--------------------------------------------------------			
--
--library IEEE;
--use IEEE.std_logic_1164.all;
--use IEEE.std_logic_arith.all;
--use IEEE.std_logic_unsigned.all;
--use IEEE.VITAL_Primitives.all;
--use IEEE.VITAL_Timing.all;
--use work.std_logic_SBT.all;
-- 
--
--entity ShiftReg427  is
-- 
--	generic ( 
--		SHIFTREG_DIV_MODE :  bit_vector(1 downto 0) := "00"  
--		);
--	port 	( 
--		clk 		: in std_logic; 
--		init 		: in std_logic; 
--		phase0 		: out std_logic; 
--		phase90		: out std_logic
--		); 
--end ShiftReg427;
--
--
--architecture  ShiftReg427_arch of ShiftReg427 is 
--
--signal ff1,ff2,ff3,ff4,ff5,ff6,ff7 : std_logic; 
--
--begin 
--
--  -- validations 	
-- initial_proc: process 
-- begin 
--  if (SHIFTREG_DIV_MODE ="10") then 
--	 assert false
--	 report "SBT_ERROR:Incorrect SHIFTREG_DIV_MODE set for simulation. The PLL Simulation results are incorrect .... " severity Error;
--   end if;
-- wait; 		-- wait forever  		
-- end process initial_proc; 
--
-- phaseshift_proc : process ( clk , init) 
-- begin 
--	if(init = '1') then 
--		ff1 <='0'; 		
--		ff2 <='0'; 		
--		ff3 <='0'; 		
--		ff4 <='1'; 		
--		ff5 <='1'; 		
--		ff6 <='1'; 		
--		ff7 <='1'; 		
--	elsif rising_edge(clk) then 
--		ff1 <= ff7; 
--	 	ff2 <= ff1;  
--		ff3 <= ff2; 
--		ff4 <= ff3;
--		if(SHIFTREG_DIV_MODE = "00" ) then 
--			ff5 <= ff4; 
--			ff6 <= ff2; 
--		elsif (SHIFTREG_DIV_MODE = "01" ) then 
--			ff5 <= ff4; 	
--			ff6 <= ff5;  
--		elsif (SHIFTREG_DIV_MODE = "11" ) then 
--			ff5 <= ff2; 
--			ff6 <= ff5; 
--	        end if ;
--		ff7 <= ff6; 
--	end if;	
-- end process  phaseshift_proc; 	
--
--	phase0 <= ff1; 	
--	phase90 <=ff2; 
--
--end ShiftReg427_arch; 

---------------------------------------------------------------------------
----			 	SbtSPLL40  				---	
---------------------------------------------------------------------------
--library IEEE;
--use IEEE.std_logic_1164.all;
--use IEEE.std_logic_arith.all;
--use IEEE.std_logic_unsigned.all;
--use IEEE.VITAL_Primitives.all;
--use IEEE.VITAL_Timing.all;
--use work.std_logic_SBT.all;
--use work.all; 
-- 
--
--entity SbtSPLL40  is
-- 
--	generic ( 
--		 FEEDBACK_PATH 			: string 		 :="SIMPLE"; 
--		 DELAY_ADJUSTMENT_MODE_FEEDBACK	: string 		 :="FIXED"; 
--		 DELAY_ADJUSTMENT_MODE_RELATIVE : string 		 :="FIXED";
--		 SHIFTREG_DIV_MODE		: bit_vector(1 downto 0) := "00"; 
--		 FDA_FEEDBACK			: bit_vector(3 downto 0) :="0000";
--		 FDA_RELATIVE			: bit_vector(3 downto 0) := "0000";
--		 PLLOUT_SELECT_PORTA		: string 		 :="GENCLK"; 
--		 PLLOUT_SELECT_PORTB            : string         	 :="GENCLK";
--
--		 DIVR				: bit_vector(3 downto 0) := "0000";
--		 DIVF  				: bit_vector(6 downto 0) := "0000000";
--		 DIVQ	   			: bit_vector(2 downto 0) := "000";  
--		 FILTER_RANGE 			: bit_vector(2 downto 0) := "000";
--		 		
-- 		 ENABLE_ICEGATE_PORTA            : bit 			 :='0';
--		 ENABLE_ICEGATE_PORTB           : bit 			 :='0' 
--	);
--	port	(
--		REFERENCECLK	: in    std_logic;
--		EXTFEEDBACK 	: in    std_logic; 				 	
--		DYNAMICDELAY	: in    std_logic_vector(7 downto 0); 
--		BYPASS 		: in	std_logic;
--		RESETB	 	: in 	std_logic;
--		PLLOUT1 	: out  	std_logic;
--		PLLOUT2		: out 	std_logic ; 
--		LOCK		: out 	std_logic  
--	); 
--
--end SbtSPLL40;
--
--	
--architecture SbtSPLL40_arch  of SbtSPLL40  is
--
--component ShiftReg427  is
-- 
--	generic ( 
--		SHIFTREG_DIV_MODE :  bit_vector(1 downto 0) := "00"  
--		);
--	port 	( 
--		clk 		: in std_logic; 
--		init 		: in std_logic; 
--		phase0 		: out std_logic; 
--		phase90		: out std_logic
--		); 
--end component;
--
--component  mux4to1   is
--	port ( 
--		a,b,c,d : in std_logic; 
--		sel 	: in std_logic_vector(1 downto 0); 
--		o	: out std_logic 
--	      ); 
--end component ;
--
--
--component FineDlyAdj  is
--	generic (
--		FIXED_DELAY_ADJUSTMENT   : bit_vector(3 downto 0) :="0000"; 
--		DELAY_ADJUSTMENT_MODE    : string 		  :="FIXED";
--		BUF_DELAY		 : time 		  := 100 ps;
--		MUXINV_DELAY		 : time 		  := 0 ps
--		); 
--	port 	( 
--		signalin		:in  std_logic; 
--		DlyAdj			:in  std_logic_vector(3 downto 0); 
--		delayedout 		:out std_logic
--		); 
--end component ;
--
-- 
--component  ABIWTCZ4  is 
--  port  	(
--                REF	:in  std_logic; 
--                FB  	:in  std_logic; 
--                FSE	:in  std_logic; 
--                BYPASS 	:in  std_logic;
--                RESET	:in  std_logic; 
--                DIVF6	:in  std_logic; 
--                DIVF5 	:in  std_logic; 
--                DIVF4 	:in  std_logic; 
--                DIVF3 	:in  std_logic; 
--                DIVF2 	:in  std_logic; 
--                DIVF1	:in  std_logic; 
--                DIVF0 	:in  std_logic; 
--                DIVQ2	:in  std_logic; 
--                DIVQ1 	:in  std_logic; 
--                DIVQ0 	:in  std_logic; 
--                DIVR3 	:in  std_logic; 
--                DIVR2 	:in  std_logic; 
--                DIVR1 	:in  std_logic; 
--                DIVR0	:in  std_logic; 
--                RANGE2  :in  std_logic; 
--                RANGE1  :in  std_logic;
--                RANGE0  :in  std_logic; 
--                LOCK    :out std_logic;
--                PLLOUT  :out std_logic  
--                );
--end component; 
--
-- signal DIVFBus    		: std_logic_vector(6 downto 0); 
-- signal DIVRBus 		: std_logic_vector(3 downto 0); 
-- signal DIVQBus 		: std_logic_vector(2 downto 0); 
-- signal RANGEBus 		: std_logic_vector(2 downto 0); 	 	
--
-- signal ABPLLOUTDiv2		: std_logic :='0'; 
-- signal ABPLLOUT     		: std_logic ; 
-- signal FSEnet       		: std_logic ; 
-- signal FBnet 	     		: std_logic ; 	
--
-- signal phase0net, phase90net  	: std_logic; 
-- signal delaymuxsel  		: std_logic_vector(1 downto 0);
-- signal pllout1Sel,pllout2Sel	: std_logic_vector(1 downto 0);	
-- signal pllout1Muxnet, pllout2Muxnet 		: std_logic; 	 
--
-- signal finedelayFBin 		: std_logic; 
-- signal finedelayFBout		: std_logic; 
-- signal fdaRelInput		: std_logic;
--
--begin 
--
-- -- generic conversions   
-- DIVFBus <= TO_STDLOGICVECTOR(DIVF); 		
-- DIVRBus <= TO_STDLOGICVECTOR(DIVR);
-- DIVQBus <= TO_STDLOGICVECTOR(DIVQ); 		
-- RANGEBus <= TO_STDLOGICVECTOR(FILTER_RANGE); 		
--  -- validations 
-- initial_proc : process 
-- begin 
-- if (PLLOUT_SELECT_PORTA = "SHIFTREG_0deg") then 
--    pllout1Sel <= "00";
-- elsif (PLLOUT_SELECT_PORTA = "SHIFTREG_90deg") then 
--    pllout1Sel <= "01";
-- elsif (PLLOUT_SELECT_PORTA = "GENCLK_HALF") then 
--    pllout1Sel <= "10";
-- elsif (PLLOUT_SELECT_PORTA = "GENCLK") then 
--    pllout1Sel <= "11";
-- else 
--        report ("************************SBT : ERROR ****************************") severity error;
--       	report ("Parameter PLLOUT_SELECT_PORTA is set to an illegal value.") severity error;
--        report ("Legal values should be one of SHIFTREG_0deg, SHIFTREG_90deg, GENCLK_HALF, GENCLK") severity error;
--        report ("Due to incorrect configuration of the PLL, the simulation results are invalid.");
-- end if ;	
--
--
--
-- if (PLLOUT_SELECT_PORTB = "SHIFTREG_0deg") then 
--    pllout2Sel <= "00";
-- elsif (PLLOUT_SELECT_PORTB = "SHIFTREG_90deg") then 
--    pllout2Sel <= "01";
-- elsif (PLLOUT_SELECT_PORTB = "GENCLK_HALF") then 
--    pllout2Sel <= "10";
-- elsif (PLLOUT_SELECT_PORTB = "GENCLK") then 
--    pllout2Sel <= "11";
-- else 
--        report ("************************SBT : ERROR ****************************") severity error;
--       	report ("Parameter PLLOUT_SELECT_PORTB is set to an illegal value.") severity error;
--        report ("Legal values should be one of SHIFTREG_0deg, SHIFTREG_90deg, GENCLK_HALF, GENCLK") severity error;
--        report ("Due to incorrect configuration of the PLL, the simulation results are invalid.");
-- end if ;	
--
--
-- -- FB 
--  if (FEEDBACK_PATH /= "EXTERNAL") then
--            report ("************************SBT : Info*****************************");
--            report ("PLL Feedback is set to INTERNAL. Any signal connected to the EXTFEEDBACK port of the PLL will be ignored");
--  end if; 
--
-- if (FEEDBACK_PATH = "EXTERNAL") then 
--       delaymuxsel <= "11";
--
--        if((DELAY_ADJUSTMENT_MODE_FEEDBACK /= "FIXED") and (DELAY_ADJUSTMENT_MODE_FEEDBACK /= "DYNAMIC") ) then 
--                report ("************************SBT : ERROR ************************");
--                report ("Since FEEDBACK_PATH=EXTERNAL, DELAY_ADJUSTMENT_MODE_FEEDBACK should be FIXED or DYNAMIC");
--                report ("Due to incorrect configuration of the PLL, the simulation results are invalid.");
--        end if; 
--        if (PLLOUT_SELECT_PORTA = "SHIFTREG_0deg" or  PLLOUT_SELECT_PORTA = "SHIFTREG_90deg" 
--			or PLLOUT_SELECT_PORTB = "SHIFTREG_0deg" or  PLLOUT_SELECT_PORTB = "SHIFTREG_90deg")  then 
--                report ("************************ SBT : ERROR **************************") severity error;
--                report ("Since FEEDBACK_PATH=EXTERNAL, Phase Adjustment is NOT permitted.") severity error;
--        end if; 
--
--   elsif (FEEDBACK_PATH = "DELAY") then 
--        delaymuxsel <= "00";
--        if ( (DELAY_ADJUSTMENT_MODE_FEEDBACK /= "FIXED") and (DELAY_ADJUSTMENT_MODE_FEEDBACK /= "DYNAMIC") ) then 
--                report ("************************ SBT : ERROR **************************") severity error ;
--                report ("Since FEEDBACK_PATH=DELAY, DELAY_ADJUSTMENT_MODE_FEEDBACK should be FIXED or DYNAMIC") severity error ;
--                report ("Due to incorrect configuration of the PLL, the simulation results are invalid.");
--        end if; 
--        if (PLLOUT_SELECT_PORTA = "SHIFTREG_0deg" or  PLLOUT_SELECT_PORTA = "SHIFTREG_90deg"
--                    or PLLOUT_SELECT_PORTB = "SHIFTREG_0deg" or PLLOUT_SELECT_PORTB = "SHIFTREG_90deg") then  
--                report ("************************ SBT : ERROR **************************") severity error;
--                report ("Since FEEDBACK_PATH=DELAY, Phase Adjustment is NOT permitted. Please set PLLOUT_SELECT_PORTA/B=GENCLK or GENCLK_HALF");
--                report ("Due to incorrect configuration of the PLL, the simulation results are invalid.");
-- 	end if;
--    elsif (FEEDBACK_PATH = "PHASE_AND_DELAY") then 
--        delaymuxsel <= "01";
--        if ( (DELAY_ADJUSTMENT_MODE_FEEDBACK /= "FIXED") and (DELAY_ADJUSTMENT_MODE_FEEDBACK /= "DYNAMIC") ) then 
--                report ("************************SBT : Attention************************");
--                report ("Since FEEDBACK_PATH=PHASE_AND_DELAY, DELAY_ADJUSTMENT_MODE_FEEDBACK should be FIXED or DYNAMIC");
--        end if; 
--        if ( (PLLOUT_SELECT_PORTA /= "SHIFTREG_0deg") and (PLLOUT_SELECT_PORTA /= "SHIFTREG_90deg" )
--                                and (PLLOUT_SELECT_PORTB /= "SHIFTREG_0deg") and  (PLLOUT_SELECT_PORTB /= "SHIFTREG_90deg") ) then 
--                report ("************************SBT : Attention************************") severity note;
--                report ("FEEDBACK_PATH=PHASE_AND_DELAY, but PLLOUT_SELECT_PORTA/B is not specified correctly") severity note;
--        end if; 
--   elsif (FEEDBACK_PATH = "SIMPLE") then 
--	-- delaymuxsel <= "00";  -- Not used 
--                -- Ignore DELAY_ADJUSTMENT_MODE_FEEDBACK, FDA_FEEDBACK
--          report ("************************SBT : Attention***************************") severity note;
--          report ("Since FEEDBACK_PATH=SIMPLE, the FDA_FEEDBACK value will be ignored") severity note;
--
--        if (PLLOUT_SELECT_PORTA = "SHIFTREG_0deg" or PLLOUT_SELECT_PORTA = "SHIFTREG_90deg"
--                   or PLLOUT_SELECT_PORTB = "SHIFTREG_0deg" or PLLOUT_SELECT_PORTB = "SHIFTREG_90deg")  then  
--                report ("************************SBT : Attention***************************") severity note;
--                report ("The PLL output frequency will be divided by 4 or 5 or 7 and phase shifted.") severity note;
--                report ("To avoid this, please set PLLOUT_SELECT_PORTA/B = GENCLK");
--        end if;
--   else
--                report ("************************SBT : Attention***************************") severity note;
--                report ("Please set FEEDBACK_PATH to a valid value. Legal settings should be one of SIMPLE, DELAY, PHASE_AND_DELAY, EXTERNAL") severity note;
--  end if; 
--
--   if( SHIFTREG_DIV_MODE ="10") then 
--                report ("************************ SBT : ERROR **************************") severity error ;
--                report ("SHIFTREG_DIV_MODE =10 is NOT permitted. Please set it 00/01/11") severity error  ;
--                report ("Due to incorrect configuration of the PLL, the simulation results are invalid.") severity error ;
--   end if; 	
-- 
-- wait ;			-- wait forever  
--
-- end process initial_proc;   
--
--  -- logic 	
--
-- ABPLLoutdiv_proc: process(ABPLLOUT) 
-- begin 
--	if rising_edge(ABPLLOUT) then 
--		ABPLLOUTDiv2 <= not(ABPLLOUTDiv2); 
--	end if ;
-- end  process ABPLLoutdiv_proc; 
--
--  -- FSE sections
-- FSEnet <= '1' when FEEDBACK_PATH = "SIMPLE" else '0';  
--
-- FBnetsel_proc:  process(finedelayFBout) 
-- begin 
--	if(FEEDBACK_PATH = "SIMPLE") then
--	   FBnet <= '0' ; 
--	else
--	   FBnet <= finedelayFBout after 1 ps;  -- 1ps delay to handle NaN  issue. 
--	end if;  	
-- end process FBnetsel_proc; 
--
--
-- instShftReg427 : ShiftReg427  
-- generic map( 
--	  	 SHIFTREG_DIV_MODE => SHIFTREG_DIV_MODE
--            )
-- port  map  (	
--                clk => ABPLLOUT, 
--                init => RESETB,
--                phase0 => phase0net, 
--                phase90 => phase90net
--            );
--
-- instFBDlyAdjInMux : mux4to1	
-- port map (
--		 a=>ABPLLOUT,
--		 b=>phase0net,
--		 c=>phase0net,
--		 d=>EXTFEEDBACK,
--		 sel=>delaymuxsel(1 downto 0),
--		 o=>finedelayFBin
--	);   
--
--
-- instPLLOUT2SelMux : mux4to1 
-- port map (
--		 a=>phase0net,
--		 b=>phase90net,
--		 c=>ABPLLOUTDiv2,
--		 d=>ABPLLOUT,
--		 sel=>pllout2Sel(1 downto 0),
--		 o=>pllout2Muxnet
--	);   
--    
-- bypasspll2_proc:  process(REFERENCECLK, pllout2Muxnet) 
-- begin 	 	
--	if(BYPASS ='1') then 
--	PLLOUT2 <= REFERENCECLK; 
--	else 
--	PLLOUT2 <= pllout2Muxnet; 
--	end if ; 
-- end process bypasspll2_proc;   
--
--	
-- instPLLOUT1SelMux : mux4to1 
-- port map (
--		 a=>phase0net,
--		 b=>phase90net,
--		 c=>ABPLLOUTDiv2,
--		 d=>ABPLLOUT,
--		 sel=>pllout1Sel(1 downto 0),
--		 o=>pllout1Muxnet
--	);   
--
--  
-- bypasspll1_proc: process(REFERENCECLK, pllout1Muxnet) 
-- begin 	 	
--	if(BYPASS ='1') then 
--	fdaRelInput <= REFERENCECLK; 
--	else 
--	fdaRelInput <= pllout1Muxnet; 
--	end if ; 
-- end process bypasspll1_proc;   
--
-- instFineDlyAdjFB : FineDlyAdj 
-- generic map    ( 
--		FIXED_DELAY_ADJUSTMENT => FDA_FEEDBACK, 
--		DELAY_ADJUSTMENT_MODE  => DELAY_ADJUSTMENT_MODE_FEEDBACK
--		)	
-- port map      (
--                DlyAdj => DYNAMICDELAY(3 downto 0),
--                signalin=>finedelayFBin,
--                delayedout=>finedelayFBout
--                );
--
-- instFineDlyAdjRel : FineDlyAdj 
-- generic map 	( 
--		FIXED_DELAY_ADJUSTMENT => FDA_RELATIVE, 
--		DELAY_ADJUSTMENT_MODE  => DELAY_ADJUSTMENT_MODE_RELATIVE
--		)		
--  port map	(
--                DlyAdj => DYNAMICDELAY(7 downto 4),
--                signalin =>fdaRelInput,
--                delayedout => PLLOUT1 
--                );
--
-- instABitsPLL : ABIWTCZ4 
-- port map  	(
--                REF => REFERENCECLK,
--                FB  => FBnet,
--                FSE => FSEnet,
--                BYPASS => BYPASS,
--                RESET => RESETB,
--                DIVF6 => DIVFBus(6),
--                DIVF5 =>DIVFBus(5),
--                DIVF4 => DIVFBus(4),
--                DIVF3 =>DIVFBus(3),
--                DIVF2 =>DIVFBus(2),
--                DIVF1 => DIVFBus(1),
--                DIVF0 => DIVFBus(0),
--                DIVQ2 => DIVQBus(2),
--                DIVQ1 => DIVQBus(1),
--                DIVQ0 => DIVQBus(0),
--                DIVR3 => DIVRBus(3),
--                DIVR2 => DIVRBus(2),
--                DIVR1 => DIVRBus(1),
--                DIVR0 => DIVRBus(0),
--                RANGE2 => RANGEBus(2),
--                RANGE1 => RANGEBus(1),
--                RANGE0 => RANGEBus(0),
--                LOCK => LOCK,
--                PLLOUT =>ABPLLOUT 
--                );
--
--end SbtSPLL40_arch;

-----------------------------------------------------------------------------------
---      		 ICE40 PLL PRIMITIVES 				   	--- 
---	#SB_PLL40_CORE	#SB_PLL40_PAD	#SB_PLL40_2_PAD	#SB_PLL40_2F_CORE   	---  		
---   	#SB_PLL40_2F_PAD	#SB_PLL40_PAD_DS   #SB_PLL40_2F_PAD_DS 	---
----------------------------------------------------------------------------------- 

---------------------------------------------------------------------------
----			 SB_PLL40_CORE	  				---	
---------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;
use work.all; 

entity SB_PLL40_CORE  is 
	
	generic ( 
		----------------------------------------------------------------------------------
                --VITAL PARAMETER
                ---------------------------------------------------------------------------------
                TimingChecksOn  	: boolean := true;
                Xon   			: boolean := true;
	        MsgOn 			: boolean := false;
                --- VITAL input port delay 
                thold_SDI_SCLK_negedge_posedge:VitalDelayType :=0 ns;
                thold_SDI_SCLK_posedge_posedge:VitalDelayType :=0 ns;
                thold_SDI_SCLK_negedge_negedge:VitalDelayType :=0 ns;
                thold_SDI_SCLK_posedge_negedge:VitalDelayType :=0 ns;
                tsetup_SDI_SCLK_negedge_posedge:VitalDelayType :=0 ns;
                tsetup_SDI_SCLK_posedge_posedge:VitalDelayType :=0 ns;
                tsetup_SDI_SCLK_negedge_negedge:VitalDelayType :=0 ns;
                tsetup_SDI_SCLK_posedge_negedge:VitalDelayType :=0 ns; 
		tpd_SCLK_SDO_negedge          	: VitalDelayType01 := (0 ns, 0 ns);				
                tipd_REFERENCECLK       : VitalDelayType01 := (0 ns, 0 ns);
            	tipd_EXTFEEDBACK        : VitalDelayType01 := (0 ns, 0 ns);
            	tipd_DYNAMICDELAY       : VitalDelayArrayType01(7 downto 0)  := (others => (0 ns, 0 ns));
            	tipd_BYPASS             : VitalDelayType01 := (0 ns, 0 ns);
            	tipd_RESETB             : VitalDelayType01 := (0 ns, 0 ns);
                tipd_SDI        	: VitalDelayType01 := (0 ns, 0 ns);
            	tipd_SCLK           	: VitalDelayType01 := (0 ns, 0 ns);
            	tipd_LATCHINPUTVALUE   	: VitalDelayType01 := (0 ns, 0 ns);
		-- VITAL Path Delay 	
            	tpd_REFERENCECLK_PLLOUTCORE           	: VitalDelayType01 := (0 ns, 0 ns);
            	tpd_REFERENCECLK_PLLOUTGLOBAL          	: VitalDelayType01 := (0 ns, 0 ns);
	         -- Entity Parameters 	
		 FEEDBACK_PATH 			: string 		 :="SIMPLE";   -- SIMPLE/DELAY/PHASE_AND_DELAY/EXTERNAL 
		 DELAY_ADJUSTMENT_MODE_FEEDBACK	: string 		 :="FIXED";    -- FIXED/DYNAMIC  
		 DELAY_ADJUSTMENT_MODE_RELATIVE : string 		 :="FIXED";    -- FIXED/DYNAMIC 
		 SHIFTREG_DIV_MODE		: bit_vector(1 downto 0) := "00";      -- 00 (div by 4)/ 01 (div by 7)/11 (div by 5)   	 
		 FDA_FEEDBACK			: bit_vector(3 downto 0) :="0000";
		 FDA_RELATIVE			: bit_vector(3 downto 0) := "0000";
		 PLLOUT_SELECT			: string 		 :="GENCLK"; 

		 DIVR				: bit_vector(3 downto 0) := "0000";
		 DIVF  				: bit_vector(6 downto 0) := "0000000";
		 DIVQ	   			: bit_vector(2 downto 0) := "000";  
		 FILTER_RANGE 			: bit_vector(2 downto 0) := "000";
		 		
 		 ENABLE_ICEGATE		        : bit 			 :='0';
		 TEST_MODE			: bit 			 :='0';  
		 EXTERNAL_DIVIDE_FACTOR         : integer 		 := 1      -- Required for PLL Config Wizard.  
	);
	port (
                REFERENCECLK		: in std_logic;           -- PLL ref clock, driven by core logic   
                PLLOUTCORE	     	: out std_logic;          -- PLL output to core logic through local routings. 
                PLLOUTGLOBAL            : out std_logic;   	  -- PLL output to dedicated global clock network
                EXTFEEDBACK             : in std_logic;  	  -- FB driven by core logic
                DYNAMICDELAY            : in std_logic_vector(7 downto 0);  -- driven by core logic
                LOCK                    : out std_logic;	  -- PLL Lock signal output  
                BYPASS                  : in std_logic; 	  -- REFCLK passed to PLLOUT when bypass is '1'.Driven by core logic
                RESETB                  : in std_logic; 	  -- Active low reset,Driven by core logic
                SDI                     : in std_logic;		  -- Test Input. Driven by core logic. 
                SDO                     : out std_logic; 	  -- Test output to RB Logic Tile.
                SCLK                    : in std_logic;	          -- Test Clk input.Driven by core logic. 
                LATCHINPUTVALUE         : in std_logic 		  -- iCEGate signal
	);

       attribute VITAL_LEVEL0 of SB_PLL40_CORE : entity is true;

end SB_PLL40_CORE; 

architecture SB_PLL40_CORE_V of SB_PLL40_CORE is 

	attribute VITAL_LEVEL0 of SB_PLL40_CORE_V  : architecture is true;


 component Sbt_DS_PLL40  is
 
	generic ( 
		 FEEDBACK_PATH 			: string 	:="SIMPLE"; 
		 DELAY_ADJUSTMENT_MODE_FEEDBACK	: string 	:="FIXED"; 
		 DELAY_ADJUSTMENT_MODE_RELATIVE : string 	:="FIXED";
		 SHIFTREG_DIV_MODE		: bit_vector(1 downto 0) := "00"; 
		 FDA_FEEDBACK			: bit_vector(3 downto 0) :="0000";
		 FDA_RELATIVE			: bit_vector(3 downto 0) := "0000";
		 PLLOUT_SELECT_PORTA		: string 	:="GENCLK"; 
		 PLLOUT_SELECT_PORTB            : string        :="GENCLK";

		 DIVR				: bit_vector(3 downto 0) := "0000";
		 DIVF  				: bit_vector(6 downto 0) := "0000000";
		 DIVQ	   			:bit_vector(2 downto 0)  := "000";  
		 FILTER_RANGE 			:bit_vector(2 downto 0)  := "000";
		 TEST_MODE         :bit        :='0'; 		
 		ENABLE_ICEGATE_PORTA             :bit 			:='0';
		ENABLE_ICEGATE_PORTB            :bit 			:='0' 
	);
	port	(
		CORE_REF_CLK	: in    std_logic;
		EXTFEEDBACK 	: in    std_logic;
		DYNAMICDELAY	: in    std_logic_vector(7 downto 0); 
		BYPASS 		: in	std_logic;
		RESETB	 	: in 	std_logic;
		PLLOUT1 	: out  	std_logic;
		PLLOUT2		: out 	std_logic ; 
		LOCK		: out 	std_logic ;
        PACKAGEPIN : in  std_logic :='0';
        PLL_SCK     :in std_logic;
        PLL_SDI     :in std_logic;
        PLL_SDO     :out std_logic 
	); 
end component;		

 component SbtSPLL40  is
 
	generic ( 
		 FEEDBACK_PATH 			: string 	:="SIMPLE"; 
		 DELAY_ADJUSTMENT_MODE_FEEDBACK	: string 	:="FIXED"; 
		 DELAY_ADJUSTMENT_MODE_RELATIVE : string 	:="FIXED";
		 SHIFTREG_DIV_MODE		: bit_vector(1 downto 0) := "00"; 
		 FDA_FEEDBACK			: bit_vector(3 downto 0) :="0000";
		 FDA_RELATIVE			: bit_vector(3 downto 0) := "0000";
		 PLLOUT_SELECT_PORTA		: string 	:="GENCLK"; 
		 PLLOUT_SELECT_PORTB            : string        :="GENCLK";

		 DIVR				: bit_vector(3 downto 0) := "0000";
		 DIVF  				: bit_vector(6 downto 0) := "0000000";
		 DIVQ	   			:bit_vector(2 downto 0)  := "000";  
		 FILTER_RANGE 			:bit_vector(2 downto 0)  := "000";
		 		
 		ENABLE_ICEGATE_PORTA             :bit 			:='0';
		ENABLE_ICEGATE_PORTB            :bit 			:='0' 
	);
	port	(
		REFERENCECLK	: in    std_logic;
		EXTFEEDBACK 	: in    std_logic;
		DYNAMICDELAY	: in    std_logic_vector(7 downto 0); 
		BYPASS 		: in	std_logic;
		RESETB	 	: in 	std_logic;
		PLLOUT1 	: out  	std_logic;
		PLLOUT2		: out 	std_logic ; 
		LOCK		: out 	std_logic  
	); 
end component;

  -- Vital Wire Delay Signals   	
  signal REFERENCECLK_ipd 	: std_ulogic := 'X';
  signal EXTFEEDBACK_ipd  	: std_ulogic := 'X';
  signal DYNAMICDELAY_ipd  	: std_logic_vector(7 downto 0) := (others =>'X');
  signal BYPASS_ipd   		: std_ulogic := 'X';
  signal RESETB_ipd 		: std_ulogic := 'X';
  signal SDI_ipd  		: std_ulogic := 'X';
  signal SCLK_ipd  		: std_ulogic := 'X';
  signal LATCHINPUTVALUE_ipd  	: std_ulogic := 'X';

 -- Vital output logic signals
 signal PLLOUTCORE_zd : std_ulogic;
 signal PLLOUTGLOBAL_zd : std_ulogic;
 signal LOCK_zd : std_ulogic;
 signal SDO_zd : std_ulogic;
 signal Violation : std_ulogic;

 -- functional signals 

 signal not_resetb  		 : std_logic; 
 signal SPLLOUT1net, SPLLOUT2net : std_logic; 
 signal PLLOUTCORE_temp 	 : std_logic; 
 signal PLLOUTGLOBAL_temp 	 : std_logic; 

begin 

 WireDelay   : block
 begin
          VitalWireDelay (REFERENCECLK_ipd, REFERENCECLK, tipd_REFERENCECLK);
          VitalWireDelay (EXTFEEDBACK_ipd,  EXTFEEDBACK, tipd_EXTFEEDBACK);
	  DYNAMIC_DELAY : for i in 7 downto 0 generate 
	          VitalWireDelay (DYNAMICDELAY_ipd(i),DYNAMICDELAY(i),tipd_DYNAMICDELAY(i));
	  end generate DYNAMIC_DELAY; 
          VitalWireDelay (BYPASS_ipd,BYPASS, tipd_BYPASS);
          VitalWireDelay (RESETB_ipd,RESETB, tipd_RESETB);
          VitalWireDelay (SDI_ipd, SDI, tipd_SDI);
          VitalWireDelay (SCLK_ipd, SCLK, tipd_SCLK);
          VitalWireDelay (LATCHINPUTVALUE_ipd, LATCHINPUTVALUE, tipd_LATCHINPUTVALUE);
 end block;

 ------ Behavioral Section   
 not_resetb <= not(RESETB_ipd);  
D: if(TEST_MODE='1') generate
 instSbtSPLL : Sbt_DS_PLL40
 generic map 	( 
		FEEDBACK_PATH 			=> FEEDBACK_PATH,
		DELAY_ADJUSTMENT_MODE_RELATIVE 	=> DELAY_ADJUSTMENT_MODE_RELATIVE,
		DELAY_ADJUSTMENT_MODE_FEEDBACK 	=> DELAY_ADJUSTMENT_MODE_FEEDBACK,
		SHIFTREG_DIV_MODE 		=> SHIFTREG_DIV_MODE,
		FDA_RELATIVE 			=> FDA_RELATIVE,
		FDA_FEEDBACK 			=> FDA_FEEDBACK,
		PLLOUT_SELECT_PORTA 		=> PLLOUT_SELECT,
		PLLOUT_SELECT_PORTB 		=> "GENCLK",
		DIVR 				=> DIVR,
		DIVF 				=> DIVF,
		DIVQ 				=> DIVQ,
		FILTER_RANGE 			=> FILTER_RANGE,
 		ENABLE_ICEGATE_PORTA             =>'0',
        	TEST_MODE          => TEST_MODE,
		ENABLE_ICEGATE_PORTB            =>'0' 
	     	)
 port map    	(
                CORE_REF_CLK 			=> REFERENCECLK_ipd,
                EXTFEEDBACK 			=> EXTFEEDBACK_ipd,
                DYNAMICDELAY 			=> DYNAMICDELAY_ipd,
                BYPASS 				=> BYPASS_ipd,
                RESETB 				=> not_resetb ,
                PLLOUT1 			=> SPLLOUT1net,
                PLLOUT2 			=> SPLLOUT2net,
                LOCK 				=> LOCK,
                PACKAGEPIN =>open,
                PLL_SCK =>      SCLK_ipd,
                PLL_SDI =>      SDI_ipd,
                PLL_SDO =>      SDO_zd
		);

end generate D;	   
S: if(TEST_MODE='0') generate
  instSbtSPLL : SbtSPLL40 
 generic map 	( 
		FEEDBACK_PATH 			=> FEEDBACK_PATH,
		DELAY_ADJUSTMENT_MODE_RELATIVE 	=> DELAY_ADJUSTMENT_MODE_RELATIVE,
		DELAY_ADJUSTMENT_MODE_FEEDBACK 	=> DELAY_ADJUSTMENT_MODE_FEEDBACK,
		SHIFTREG_DIV_MODE 		=> SHIFTREG_DIV_MODE,
		FDA_RELATIVE 			=> FDA_RELATIVE,
		FDA_FEEDBACK 			=> FDA_FEEDBACK,
		PLLOUT_SELECT_PORTA 		=> PLLOUT_SELECT,
		PLLOUT_SELECT_PORTB 		=> "GENCLK",
		DIVR 				=> DIVR,
		DIVF 				=> DIVF,
		DIVQ 				=> DIVQ,
		FILTER_RANGE 			=> FILTER_RANGE,
 		ENABLE_ICEGATE_PORTA            =>'0',		
		ENABLE_ICEGATE_PORTB            =>'0' 
	     	)
 port map    	(
                REFERENCECLK 			=> REFERENCECLK_ipd,
                EXTFEEDBACK 			=> EXTFEEDBACK_ipd,
                DYNAMICDELAY 			=> DYNAMICDELAY_ipd,
                BYPASS 				=> BYPASS_ipd,
                RESETB 				=> not_resetb ,
                PLLOUT1 			=> SPLLOUT1net,
                PLLOUT2 			=> SPLLOUT2net,
                LOCK 				=> LOCK
		);


end generate S;

 process(PLLOUTCORE_temp, SPLLOUT1net)  
 begin 
	if(ENABLE_ICEGATE = '1' and LATCHINPUTVALUE_ipd ='1') then 
		PLLOUTCORE_temp <= PLLOUTCORE_temp ; 
	else 
		PLLOUTCORE_temp <= SPLLOUT1net; 
	end if;
 end process; 


 process(PLLOUTGLOBAL_temp, SPLLOUT1net)  
 begin 
	if(ENABLE_ICEGATE = '1' and LATCHINPUTVALUE_ipd ='1') then 
		PLLOUTGLOBAL_temp <= PLLOUTGLOBAL_temp ; 
	else 
		PLLOUTGLOBAL_temp <= SPLLOUT1net; 
	end if; 
 end process; 

 PLLOUTCORE_zd 	<= PLLOUTCORE_temp; 
 PLLOUTGLOBAL_zd 	<= PLLOUTGLOBAL_temp;  

 
 ---------------------------- 
 -- Vital Path delay  
 ---------------------------
 VITALTimingCheck:process(SCLK_ipd,SDI_ipd)
     variable Tviol_SDI_SCLK_posedge       	: std_ulogic := '0';
     variable Tmkr_SDI_SCLK_posedge       	: VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_SDI_SCLK_negedge       	: std_ulogic := '0';
     variable Tmkr_SDI_SCLK_negedge       	: VitalTimingDataType := VitalTimingDataInit;
 begin
 if(TimingChecksOn) then
           VitalSetupHoldCheck (
        Violation      => Tviol_SDI_SCLK_posedge,
        TimingData     => Tmkr_SDI_SCLK_posedge,
        TestSignal     => SDI_ipd,
        TestSignalName => "SDI",
        TestDelay      => 0 ns,
        RefSignal      => SCLK_ipd,
        RefSignalName  => "SCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_SDI_SCLK_posedge_posedge,
        SetupLow       => tsetup_SDI_SCLK_negedge_posedge,
        HoldLow        => thold_SDI_SCLK_posedge_posedge,
        HoldHigh       => thold_SDI_SCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/PLL40",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

           VitalSetupHoldCheck (
        Violation      => Tviol_SDI_SCLK_negedge,
        TimingData     => Tmkr_SDI_SCLK_negedge,
        TestSignal     => SDI_ipd,
        TestSignalName => "SDI",
        TestDelay      => 0 ns,
        RefSignal      => SCLK_ipd,
        RefSignalName  => "SCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_SDI_SCLK_posedge_negedge,
        SetupLow       => tsetup_SDI_SCLK_negedge_negedge,
        HoldLow        => thold_SDI_SCLK_posedge_negedge,
        HoldHigh       => thold_SDI_SCLK_negedge_negedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/PLL40",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
end if;
end process VITALTimingCheck;

  VITALPathDelay          : process (PLLOUTCORE_zd, PLLOUTGLOBAL_zd, REFERENCECLK_ipd,SCLK_ipd,SDO_zd )
  	variable PLLOUTCORE_GlitchData 	 : VitalGlitchDataType;
	variable PLLOUTCORE_sig : std_ulogic := 'X';
	variable PLLOUTGLOBAL_GlitchData : VitalGlitchDataType;
	variable PLLOUTGLOBAL_sig : std_ulogic := 'X';
	variable SDO_GlitchData : VitalGlitchDataType;
	variable SDO_sig : std_ulogic := 'X';
	variable LOCK_zd		 : VitalGlitchDataType;

  begin 		
  PLLOUTCORE_sig:=PLLOUTCORE_zd;
  PLLOUTGLOBAL_sig:=PLLOUTGLOBAL_zd;
  SDO_sig:=SDO_zd;
  VitalPathDelay01 (
      OutSignal                 => PLLOUTCORE,
      GlitchData                => PLLOUTCORE_GlitchData,
      OutSignalName             => "PLLOUTCORE",
      OutTemp                   => PLLOUTCORE_sig,
      Paths                     => (0 => (REFERENCECLK_ipd'last_event, tpd_REFERENCECLK_PLLOUTCORE,true)
							),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
	  
      VitalPathDelay01 (
      OutSignal                 => PLLOUTGLOBAL,
      GlitchData                => PLLOUTGLOBAL_GlitchData,
      OutSignalName             => "PLLOUTGLOBAL",
      OutTemp                   => PLLOUTGLOBAL_sig,
      Paths                     => (0 => (REFERENCECLK_ipd'last_event, tpd_REFERENCECLK_PLLOUTGLOBAL, true)
									),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
	  
	        VitalPathDelay01 (
      OutSignal                 => SDO,
      GlitchData                => SDO_GlitchData,
      OutSignalName             => "SDO",
      OutTemp                   => SDO_sig,
      Paths                     => (0 => (SCLK_ipd'last_event, tpd_SCLK_SDO_negedge, true)
									),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
 end process VITALPathDelay;	

end SB_PLL40_CORE_V; 



---------------------------------------------------------------------------
----			 SB_PLL40_PAD	  				---	
---------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;
use work.all; 

entity SB_PLL40_PAD  is 
	
	generic ( 
		----------------------------------------------------------------------------------
                --VITAL PARAMETER
                ---------------------------------------------------------------------------------
                TimingChecksOn  	: boolean := true;
                Xon   			: boolean := true;
	        MsgOn 			: boolean := false;
			--- VITAL input port delay 		   
                thold_SDI_SCLK_negedge_posedge:VitalDelayType :=0 ns;
                thold_SDI_SCLK_posedge_posedge:VitalDelayType :=0 ns;
                thold_SDI_SCLK_negedge_negedge:VitalDelayType :=0 ns;
                thold_SDI_SCLK_posedge_negedge:VitalDelayType :=0 ns;
                tsetup_SDI_SCLK_negedge_posedge:VitalDelayType :=0 ns;
                tsetup_SDI_SCLK_posedge_posedge:VitalDelayType :=0 ns;
                tsetup_SDI_SCLK_negedge_negedge:VitalDelayType :=0 ns;
                tsetup_SDI_SCLK_posedge_negedge:VitalDelayType :=0 ns; 
				tpd_SCLK_SDO_negedge          	: VitalDelayType01 := (0 ns, 0 ns);				
                tipd_PACKAGEPIN       : VitalDelayType01 := (0 ns, 0 ns);
            	tipd_EXTFEEDBACK        : VitalDelayType01 := (0 ns, 0 ns);
            	tipd_DYNAMICDELAY       : VitalDelayArrayType01(7 downto 0)  := (others => (0 ns, 0 ns));
            	tipd_BYPASS             : VitalDelayType01 := (0 ns, 0 ns);
            	tipd_RESETB             : VitalDelayType01 := (0 ns, 0 ns);
                tipd_SDI        	: VitalDelayType01 := (0 ns, 0 ns);
            	tipd_SCLK           	: VitalDelayType01 := (0 ns, 0 ns);
            	tipd_LATCHINPUTVALUE   	: VitalDelayType01 := (0 ns, 0 ns);
		-- VITAL Path Delay 	
            	tpd_PACKAGEPIN_PLLOUTCORE           	: VitalDelayType01 := (0 ns, 0 ns);
            	tpd_PACKAGEPIN_PLLOUTGLOBAL          	: VitalDelayType01 := (0 ns, 0 ns);
	         -- Entity Parameters 	
		 FEEDBACK_PATH 			: string 		 :="SIMPLE";   -- SIMPLE/DELAY/PHASE_AND_DELAY/EXTERNAL 
		 DELAY_ADJUSTMENT_MODE_FEEDBACK	: string 		 :="FIXED";    -- FIXED/DYNAMIC  
		 DELAY_ADJUSTMENT_MODE_RELATIVE : string 		 :="FIXED";    -- FIXED/DYNAMIC 
		 SHIFTREG_DIV_MODE		: bit_vector(1 downto 0) := "00";      -- 00 (div by 4)/ 01 (div by 7)/11 (div by 5)   	 
		 FDA_FEEDBACK			: bit_vector(3 downto 0) :="0000";
		 FDA_RELATIVE			: bit_vector(3 downto 0) := "0000";
		 PLLOUT_SELECT			: string 		 :="GENCLK"; 

		 DIVR				: bit_vector(3 downto 0) := "0000";
		 DIVF  				: bit_vector(6 downto 0) := "0000000";
		 DIVQ	   			: bit_vector(2 downto 0) := "000";  
		 FILTER_RANGE 			: bit_vector(2 downto 0) := "000";
		 		
 		 ENABLE_ICEGATE		        : bit 			 :='0';
		 TEST_MODE			: bit 			 :='0';  
		 EXTERNAL_DIVIDE_FACTOR         : integer 		 := 1      -- Required for PLL Config Wizard.  
	);
	port (
                PACKAGEPIN		: in std_logic;           -- PLL ref clock, driven by PAD.  
                PLLOUTCORE	     	: out std_logic;          -- PLL output to core logic through local routings. 
                PLLOUTGLOBAL            : out std_logic;   	  -- PLL output to dedicated global clock network
                EXTFEEDBACK             : in std_logic;  	  -- FB driven by core logic
                DYNAMICDELAY            : in std_logic_vector(7 downto 0);  -- driven by core logic
                LOCK                    : out std_logic;	  -- PLL Lock signal output  
                BYPASS                  : in std_logic; 	  -- REFCLK passed to PLLOUT when bypass is '1'.Driven by core logic
                RESETB                  : in std_logic; 	  -- Active low reset,Driven by core logic
                SDI                     : in std_logic;		  -- Test Input. Driven by core logic. 
                SDO                     : out std_logic; 	  -- Test output to RB Logic Tile.
                SCLK                    : in std_logic;	          -- Test Clk input.Driven by core logic. 
                LATCHINPUTVALUE         : in std_logic 		  -- iCEGate signal
	);

       attribute VITAL_LEVEL0 of SB_PLL40_PAD : entity is true;

end SB_PLL40_PAD; 

architecture SB_PLL40_PAD_V of SB_PLL40_PAD is 

	attribute VITAL_LEVEL0 of SB_PLL40_PAD_V  : architecture is true;

 component Sbt_DS_PLL40  is
 
	generic ( 
		 FEEDBACK_PATH 			: string 	:="SIMPLE"; 
		 DELAY_ADJUSTMENT_MODE_FEEDBACK	: string 	:="FIXED"; 
		 DELAY_ADJUSTMENT_MODE_RELATIVE : string 	:="FIXED";
		 SHIFTREG_DIV_MODE		: bit_vector(1 downto 0) := "00"; 
		 FDA_FEEDBACK			: bit_vector(3 downto 0) :="0000";
		 FDA_RELATIVE			: bit_vector(3 downto 0) := "0000";
		 PLLOUT_SELECT_PORTA		: string 	:="GENCLK"; 
		 PLLOUT_SELECT_PORTB            : string        :="GENCLK";

		 DIVR				: bit_vector(3 downto 0) := "0000";
		 DIVF  				: bit_vector(6 downto 0) := "0000000";
		 DIVQ	   			:bit_vector(2 downto 0)  := "000";  
		 FILTER_RANGE 			:bit_vector(2 downto 0)  := "000";
		 TEST_MODE         :bit        :='0'; 		
 		ENABLE_ICEGATE_PORTA             :bit 			:='0';
		ENABLE_ICEGATE_PORTB            :bit 			:='0' 
	);
	port	(
		CORE_REF_CLK	: in    std_logic:='0';
		EXTFEEDBACK 	: in    std_logic;
		DYNAMICDELAY	: in    std_logic_vector(7 downto 0); 
		BYPASS 		: in	std_logic;
		RESETB	 	: in 	std_logic;
		PLLOUT1 	: out  	std_logic;
		PLLOUT2		: out 	std_logic ; 
		LOCK		: out 	std_logic ;
        PACKAGEPIN : in  std_logic :='0';
        PLL_SCK     :in std_logic;
        PLL_SDI     :in std_logic;
        PLL_SDO     :out std_logic 
	); 
end component;	
 component SbtSPLL40  is
 
	generic ( 
		 FEEDBACK_PATH 			: string 	:="SIMPLE"; 
		 DELAY_ADJUSTMENT_MODE_FEEDBACK	: string 	:="FIXED"; 
		 DELAY_ADJUSTMENT_MODE_RELATIVE : string 	:="FIXED";
		 SHIFTREG_DIV_MODE		: bit_vector(1 downto 0) := "00"; 
		 FDA_FEEDBACK			: bit_vector(3 downto 0) :="0000";
		 FDA_RELATIVE			: bit_vector(3 downto 0) := "0000";
		 PLLOUT_SELECT_PORTA		: string 	:="GENCLK"; 
		 PLLOUT_SELECT_PORTB            : string        :="GENCLK";

		 DIVR				: bit_vector(3 downto 0) := "0000";
		 DIVF  				: bit_vector(6 downto 0) := "0000000";
		 DIVQ	   			:bit_vector(2 downto 0)  := "000";  
		 FILTER_RANGE 			:bit_vector(2 downto 0)  := "000";
		 		
 		ENABLE_ICEGATE_PORTA             :bit 			:='0';
		ENABLE_ICEGATE_PORTB            :bit 			:='0' 
	);
	port	(
		REFERENCECLK	: in    std_logic;
		EXTFEEDBACK 	: in    std_logic;
		DYNAMICDELAY	: in    std_logic_vector(7 downto 0); 
		BYPASS 		: in	std_logic;
		RESETB	 	: in 	std_logic;
		PLLOUT1 	: out  	std_logic;
		PLLOUT2		: out 	std_logic ; 
		LOCK		: out 	std_logic  
	); 
end component;

  -- Vital Wire Delay Signals   	
  signal PACKAGEPIN_ipd 	: std_ulogic := 'X';
  signal EXTFEEDBACK_ipd  	: std_ulogic := 'X';
  signal DYNAMICDELAY_ipd  	: std_logic_vector(7 downto 0) := (others =>'X');
  signal BYPASS_ipd   		: std_ulogic := 'X';
  signal RESETB_ipd 		: std_ulogic := 'X';
  signal SDI_ipd  		: std_ulogic := 'X';
  signal SCLK_ipd  		: std_ulogic := 'X';
  signal LATCHINPUTVALUE_ipd  	: std_ulogic := 'X';

 -- Vital output logic signals
 signal PLLOUTCORE_zd : std_ulogic;
 signal PLLOUTGLOBAL_zd : std_ulogic;
 signal LOCK_zd : std_ulogic;
 signal SDO_zd : std_ulogic;
 signal Violation : std_ulogic;

 -- Functional Signals 
 signal not_resetb  		 : std_logic; 
 signal SPLLOUT1net, SPLLOUT2net : std_logic; 
 signal PLLOUTCORE_temp 	 : std_logic; 
 signal PLLOUTGLOBAL_temp 	 : std_logic; 

begin 

 WireDelay   : block
 begin
          VitalWireDelay (PACKAGEPIN_ipd, PACKAGEPIN, tipd_PACKAGEPIN);
          VitalWireDelay (EXTFEEDBACK_ipd,  EXTFEEDBACK, tipd_EXTFEEDBACK);
	  DYNAMIC_DELAY : for i in 7 downto 0 generate 
	          VitalWireDelay (DYNAMICDELAY_ipd(i),DYNAMICDELAY(i),tipd_DYNAMICDELAY(i));
	  end generate DYNAMIC_DELAY; 
          VitalWireDelay (BYPASS_ipd,BYPASS, tipd_BYPASS);
          VitalWireDelay (RESETB_ipd,RESETB, tipd_RESETB);
          VitalWireDelay (SDI_ipd, SDI, tipd_SDI);
          VitalWireDelay (SCLK_ipd, SCLK, tipd_SCLK);
          VitalWireDelay (LATCHINPUTVALUE_ipd, LATCHINPUTVALUE, tipd_LATCHINPUTVALUE);
 end block;

 ------ Behavioral Section   
 not_resetb <= not(RESETB_ipd);  
 D: if(TEST_MODE='1') generate
 instSbtSPLL : Sbt_DS_PLL40
 generic map 	( 
		FEEDBACK_PATH 			=> FEEDBACK_PATH,
		DELAY_ADJUSTMENT_MODE_RELATIVE 	=> DELAY_ADJUSTMENT_MODE_RELATIVE,
		DELAY_ADJUSTMENT_MODE_FEEDBACK 	=> DELAY_ADJUSTMENT_MODE_FEEDBACK,
		SHIFTREG_DIV_MODE 		=> SHIFTREG_DIV_MODE,
		FDA_RELATIVE 			=> FDA_RELATIVE,
		FDA_FEEDBACK 			=> FDA_FEEDBACK,
		PLLOUT_SELECT_PORTA 		=> PLLOUT_SELECT,
		PLLOUT_SELECT_PORTB 		=> "GENCLK",
		DIVR 				=> DIVR,
		DIVF 				=> DIVF,
		DIVQ 				=> DIVQ,
		FILTER_RANGE 			=> FILTER_RANGE,
 		ENABLE_ICEGATE_PORTA             =>'0',
        	TEST_MODE          => TEST_MODE,
		ENABLE_ICEGATE_PORTB            =>'0' 
	     	)
 port map    	(
                CORE_REF_CLK 			=>open,
                EXTFEEDBACK 			=> EXTFEEDBACK_ipd,
                DYNAMICDELAY 			=> DYNAMICDELAY_ipd,
                BYPASS 				=> BYPASS_ipd,
                RESETB 				=> not_resetb ,
                PLLOUT1 			=> SPLLOUT1net,
                PLLOUT2 			=> SPLLOUT2net,
                LOCK 				=> LOCK,
                PACKAGEPIN =>PACKAGEPIN_ipd,
                PLL_SCK =>      SCLK_ipd,
                PLL_SDI =>      SDI_ipd,
                PLL_SDO =>      SDO_zd
		);
end generate D;	
S: if(TEST_MODE='0') generate
 instSbtSPLL : SbtSPLL40 
 generic map 	( 
		FEEDBACK_PATH 			=> FEEDBACK_PATH,
		DELAY_ADJUSTMENT_MODE_RELATIVE 	=> DELAY_ADJUSTMENT_MODE_RELATIVE,
		DELAY_ADJUSTMENT_MODE_FEEDBACK 	=> DELAY_ADJUSTMENT_MODE_FEEDBACK,
		SHIFTREG_DIV_MODE 		=> SHIFTREG_DIV_MODE,
		FDA_RELATIVE 			=> FDA_RELATIVE,
		FDA_FEEDBACK 			=> FDA_FEEDBACK,
		PLLOUT_SELECT_PORTA 		=> PLLOUT_SELECT,
		PLLOUT_SELECT_PORTB 		=> "GENCLK",
		DIVR 				=> DIVR,
		DIVF 				=> DIVF,
		DIVQ 				=> DIVQ,
		FILTER_RANGE 			=> FILTER_RANGE,
 		ENABLE_ICEGATE_PORTA            =>'0',
		ENABLE_ICEGATE_PORTB            =>'0' 
	     	)
 port map    	(
                REFERENCECLK 			=> PACKAGEPIN_ipd,
                EXTFEEDBACK 			=> EXTFEEDBACK_ipd,
                DYNAMICDELAY 			=> DYNAMICDELAY_ipd,
                BYPASS 				=> BYPASS_ipd,
                RESETB 				=> not_resetb ,
                PLLOUT1 			=> SPLLOUT1net,
                PLLOUT2 			=> SPLLOUT2net,
                LOCK 				=> LOCK
		);
 end generate S;	


 process(PLLOUTCORE_temp, SPLLOUT1net)  
 begin 
	if(ENABLE_ICEGATE = '1' and LATCHINPUTVALUE_ipd ='1') then 
		PLLOUTCORE_temp <= PLLOUTCORE_temp ; 
	else 
		PLLOUTCORE_temp <= SPLLOUT1net; 
	end if;
 end process; 


 process(PLLOUTGLOBAL_temp, SPLLOUT1net)  
 begin 
	if(ENABLE_ICEGATE = '1' and LATCHINPUTVALUE_ipd ='1') then 
		PLLOUTGLOBAL_temp <= PLLOUTGLOBAL_temp ; 
	else 
		PLLOUTGLOBAL_temp <= SPLLOUT1net; 
	end if; 
 end process; 

 PLLOUTCORE_zd 	<= PLLOUTCORE_temp; 
 PLLOUTGLOBAL_zd 	<= PLLOUTGLOBAL_temp;  

 VITALTimingCheck:process(SCLK_ipd,SDI_ipd)
     variable Tviol_SDI_SCLK_posedge       	: std_ulogic := '0';
     variable Tmkr_SDI_SCLK_posedge       	: VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_SDI_SCLK_negedge       	: std_ulogic := '0';
     variable Tmkr_SDI_SCLK_negedge       	: VitalTimingDataType := VitalTimingDataInit;
 begin
 if(TimingChecksOn) then
           VitalSetupHoldCheck (
        Violation      => Tviol_SDI_SCLK_posedge,
        TimingData     => Tmkr_SDI_SCLK_posedge,
        TestSignal     => SDI_ipd,
        TestSignalName => "SDI",
        TestDelay      => 0 ns,
        RefSignal      => SCLK_ipd,
        RefSignalName  => "SCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_SDI_SCLK_posedge_posedge,
        SetupLow       => tsetup_SDI_SCLK_negedge_posedge,
        HoldLow        => thold_SDI_SCLK_posedge_posedge,
        HoldHigh       => thold_SDI_SCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/PLL40",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

           VitalSetupHoldCheck (
        Violation      => Tviol_SDI_SCLK_negedge,
        TimingData     => Tmkr_SDI_SCLK_negedge,
        TestSignal     => SDI_ipd,
        TestSignalName => "SDI",
        TestDelay      => 0 ns,
        RefSignal      => SCLK_ipd,
        RefSignalName  => "SCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_SDI_SCLK_posedge_negedge,
        SetupLow       => tsetup_SDI_SCLK_negedge_negedge,
        HoldLow        => thold_SDI_SCLK_posedge_negedge,
        HoldHigh       => thold_SDI_SCLK_negedge_negedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/PLL40",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
end if;
end process VITALTimingCheck; 
 ---------------------------- 
 -- Vital Path delay  
 ---------------------------
  VITALPathDelay          : process (PLLOUTCORE_zd, PLLOUTGLOBAL_zd, PACKAGEPIN_ipd,SCLK_ipd,SDO_zd )
  	variable PLLOUTCORE_GlitchData 	 : VitalGlitchDataType;
	variable PLLOUTCORE_sig : std_ulogic := 'X';
	variable PLLOUTGLOBAL_GlitchData : VitalGlitchDataType;
	variable PLLOUTGLOBAL_sig : std_ulogic := 'X';
	variable SDO_GlitchData : VitalGlitchDataType;
	variable SDO_sig : std_ulogic := 'X';
	variable LOCK_zd		 : VitalGlitchDataType;

  begin 	
	  PLLOUTCORE_sig:=PLLOUTCORE_zd;
  PLLOUTGLOBAL_sig:=PLLOUTGLOBAL_zd;
  SDO_sig:=SDO_zd;
  VitalPathDelay01 (
      OutSignal                 => PLLOUTCORE,
      GlitchData                => PLLOUTCORE_GlitchData,
      OutSignalName             => "PLLOUTCORE",
      OutTemp                   => PLLOUTCORE_sig,
      Paths                     => (0 => (PACKAGEPIN_ipd'last_event, tpd_PACKAGEPIN_PLLOUTCORE,true)
							),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
	  
      VitalPathDelay01 (
      OutSignal                 => PLLOUTGLOBAL,
      GlitchData                => PLLOUTGLOBAL_GlitchData,
      OutSignalName             => "PLLOUTGLOBAL",
      OutTemp                   => PLLOUTGLOBAL_sig,
      Paths                     => (0 => (PACKAGEPIN_ipd'last_event, tpd_PACKAGEPIN_PLLOUTGLOBAL, true)
									),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
	        VitalPathDelay01 (
      OutSignal                 => SDO,
      GlitchData                => SDO_GlitchData,
      OutSignalName             => "SDO",
      OutTemp                   => SDO_sig,
      Paths                     => (0 => (SCLK_ipd'last_event, tpd_SCLK_SDO_negedge, true)
									),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
  end process VITALPathDelay;	

end SB_PLL40_PAD_V; 
 


---------------------------------------------------------------------------
----			 SB_PLL40_2_PAD	  				---	
---------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;
use work.all; 

entity SB_PLL40_2_PAD  is 
	
	generic ( 
		----------------------------------------------------------------------------------
                --VITAL PARAMETER
                ---------------------------------------------------------------------------------
                TimingChecksOn  	: boolean := true;
                Xon   			: boolean := true;
	        MsgOn 			: boolean := false;	 
                thold_SDI_SCLK_negedge_posedge:VitalDelayType :=0 ns;
                thold_SDI_SCLK_posedge_posedge:VitalDelayType :=0 ns;
                thold_SDI_SCLK_negedge_negedge:VitalDelayType :=0 ns;
                thold_SDI_SCLK_posedge_negedge:VitalDelayType :=0 ns;
                tsetup_SDI_SCLK_negedge_posedge:VitalDelayType :=0 ns;
                tsetup_SDI_SCLK_posedge_posedge:VitalDelayType :=0 ns;
                tsetup_SDI_SCLK_negedge_negedge:VitalDelayType :=0 ns;
                tsetup_SDI_SCLK_posedge_negedge:VitalDelayType :=0 ns; 
				tpd_SCLK_SDO_negedge          	: VitalDelayType01 := (0 ns, 0 ns);	
                --- VITAL input port delay 
                tipd_PACKAGEPIN       : VitalDelayType01 := (0 ns, 0 ns);
            	tipd_EXTFEEDBACK        : VitalDelayType01 := (0 ns, 0 ns);
            	tipd_DYNAMICDELAY       : VitalDelayArrayType01(7 downto 0)  := (others => (0 ns, 0 ns));
            	tipd_BYPASS             : VitalDelayType01 := (0 ns, 0 ns);
            	tipd_RESETB             : VitalDelayType01 := (0 ns, 0 ns);
                tipd_SDI        	: VitalDelayType01 := (0 ns, 0 ns);
            	tipd_SCLK           	: VitalDelayType01 := (0 ns, 0 ns);
            	tipd_LATCHINPUTVALUE   	: VitalDelayType01 := (0 ns, 0 ns);
		-- VITAL Path Delay 	
            	tpd_PACKAGEPIN_PLLOUTCOREA           	: VitalDelayType01 := (0 ns, 0 ns);
            	tpd_PACKAGEPIN_PLLOUTGLOBALA          	: VitalDelayType01 := (0 ns, 0 ns);

            	tpd_PACKAGEPIN_PLLOUTCOREB           	: VitalDelayType01 := (0 ns, 0 ns);
            	tpd_PACKAGEPIN_PLLOUTGLOBALB          	: VitalDelayType01 := (0 ns, 0 ns);
	         -- Entity Parameters 	
		 FEEDBACK_PATH 			: string 		 :="SIMPLE";   -- SIMPLE/DELAY/PHASE_AND_DELAY/EXTERNAL 
		 DELAY_ADJUSTMENT_MODE_FEEDBACK	: string 		 :="FIXED";    -- FIXED/DYNAMIC  
		 DELAY_ADJUSTMENT_MODE_RELATIVE : string 		 :="FIXED";    -- FIXED/DYNAMIC 
		 SHIFTREG_DIV_MODE		: bit_vector(1 downto 0) := "00";      -- 00 (div by 4)/ 01 (div by 7)/11 (div by 5)   	 
		 FDA_FEEDBACK			: bit_vector(3 downto 0) :="0000";
		 FDA_RELATIVE			: bit_vector(3 downto 0) := "0000";
		 PLLOUT_SELECT_PORTB		: string 		 :="GENCLK"; 

		 DIVR				: bit_vector(3 downto 0) := "0000";
		 DIVF  				: bit_vector(6 downto 0) := "0000000";
		 DIVQ	   			: bit_vector(2 downto 0) := "000";  
		 FILTER_RANGE 			: bit_vector(2 downto 0) := "000";
		 		
 		 ENABLE_ICEGATE_PORTA	        : bit 			 :='0';
 		 ENABLE_ICEGATE_PORTB	        : bit 			 :='0';
		 TEST_MODE			: bit 			 :='0';  
		 EXTERNAL_DIVIDE_FACTOR         : integer 		 := 1      -- Required for PLL Config Wizard.  
	);
	port (
                PACKAGEPIN		: in std_logic;           -- PLL ref clock, driven by PAD.  
                PLLOUTCOREA	     	: out std_logic;          -- PLLA output to core logic through local routings. 
                PLLOUTGLOBALA           : out std_logic;   	  -- PLLA output to dedicated global clock network
                PLLOUTCOREB	     	: out std_logic;          -- PLLB output to core logic through local routings. 
                PLLOUTGLOBALB           : out std_logic;   	  -- PLLB output to dedicated global clock network
                EXTFEEDBACK             : in std_logic;  	  -- FB driven by core logic
                DYNAMICDELAY            : in std_logic_vector(7 downto 0);  -- driven by core logic
                LOCK                    : out std_logic;	  -- PLL Lock signal output  
                BYPASS                  : in std_logic; 	  -- REFCLK passed to PLLOUT when bypass is '1'.Driven by core logic
                RESETB                  : in std_logic; 	  -- Active low reset,Driven by core logic
                SDI                     : in std_logic;		  -- Test Input. Driven by core logic. 
                SDO                     : out std_logic; 	  -- Test output to RB Logic Tile.
                SCLK                    : in std_logic;	          -- Test Clk input.Driven by core logic. 
                LATCHINPUTVALUE         : in std_logic 		  -- iCEGate signal
	);

       attribute VITAL_LEVEL0 of SB_PLL40_2_PAD : entity is true;

end SB_PLL40_2_PAD; 

architecture SB_PLL40_2_PAD_V of SB_PLL40_2_PAD is 

	attribute VITAL_LEVEL0 of SB_PLL40_2_PAD_V  : architecture is true;


 component SbtSPLL40  is
 
	generic ( 
		 FEEDBACK_PATH 			: string 	:="SIMPLE"; 
		 DELAY_ADJUSTMENT_MODE_FEEDBACK	: string 	:="FIXED"; 
		 DELAY_ADJUSTMENT_MODE_RELATIVE : string 	:="FIXED";
		 SHIFTREG_DIV_MODE		: bit_vector(1 downto 0) := "00";		 
		 FDA_FEEDBACK			: bit_vector(3 downto 0) :="0000";
		 FDA_RELATIVE			: bit_vector(3 downto 0) := "0000";
		 PLLOUT_SELECT_PORTA		: string 	:="GENCLK"; 
		 PLLOUT_SELECT_PORTB            : string        :="GENCLK"; 

		 DIVR				: bit_vector(3 downto 0) := "0000";
		 DIVF  				: bit_vector(6 downto 0) := "0000000";
		 DIVQ	   			:bit_vector(2 downto 0)  := "000";  
		 FILTER_RANGE 			:bit_vector(2 downto 0)  := "000";
		 		
 		ENABLE_ICEGATE_PORTA             :bit 			:='0';
		ENABLE_ICEGATE_PORTB            :bit 			:='0' 
	);
	port	(
		REFERENCECLK	: in    std_logic;
		EXTFEEDBACK 	: in    std_logic;
		DYNAMICDELAY	: in    std_logic_vector(7 downto 0); 
		BYPASS 		: in	std_logic;
		RESETB	 	: in 	std_logic;
		PLLOUT1 	: out  	std_logic;
		PLLOUT2		: out 	std_logic ; 
		LOCK		: out 	std_logic  
	); 
end component;

component Sbt_DS_PLL40  is
 
	generic ( 
		 FEEDBACK_PATH 			: string 	:="SIMPLE"; 
		 DELAY_ADJUSTMENT_MODE_FEEDBACK	: string 	:="FIXED"; 
		 DELAY_ADJUSTMENT_MODE_RELATIVE : string 	:="FIXED";
		 SHIFTREG_DIV_MODE		: bit_vector(1 downto 0) := "00"; 
		 FDA_FEEDBACK			: bit_vector(3 downto 0) :="0000";
		 FDA_RELATIVE			: bit_vector(3 downto 0) := "0000";
		 PLLOUT_SELECT_PORTA		: string 	:="GENCLK"; 
		 PLLOUT_SELECT_PORTB            : string        :="GENCLK";

		 DIVR				: bit_vector(3 downto 0) := "0000";
		 DIVF  				: bit_vector(6 downto 0) := "0000000";
		 DIVQ	   			:bit_vector(2 downto 0)  := "000";  
		 FILTER_RANGE 			:bit_vector(2 downto 0)  := "000";
		 TEST_MODE         :bit        :='0'; 		
 		ENABLE_ICEGATE_PORTA             :bit 			:='0';
		ENABLE_ICEGATE_PORTB            :bit 			:='0' 
	);
	port	(
		CORE_REF_CLK	: in    std_logic:='0';
		EXTFEEDBACK 	: in    std_logic;
		DYNAMICDELAY	: in    std_logic_vector(7 downto 0); 
		BYPASS 		: in	std_logic;
		RESETB	 	: in 	std_logic;
		PLLOUT1 	: out  	std_logic;
		PLLOUT2		: out 	std_logic ; 
		LOCK		: out 	std_logic ;
        PACKAGEPIN : in  std_logic :='0';
        PLL_SCK     :in std_logic;
        PLL_SDI     :in std_logic;
        PLL_SDO     :out std_logic 
	); 
end component;	
  -- Vital Wire Delay Signals   	
  signal PACKAGEPIN_ipd 	: std_ulogic := 'X';
  signal EXTFEEDBACK_ipd  	: std_ulogic := 'X';
  signal DYNAMICDELAY_ipd  	: std_logic_vector(7 downto 0) := (others =>'X');
  signal BYPASS_ipd   		: std_ulogic := 'X';
  signal RESETB_ipd 		: std_ulogic := 'X';
  signal SDI_ipd  		: std_ulogic := 'X';
  signal SCLK_ipd  		: std_ulogic := 'X';
  signal LATCHINPUTVALUE_ipd  	: std_ulogic := 'X';

 -- Vital output logic signals
 signal PLLOUTCOREA_zd : std_ulogic;
 signal PLLOUTGLOBALA_zd : std_ulogic;
 signal PLLOUTCOREB_zd : std_ulogic;
 signal PLLOUTGLOBALB_zd : std_ulogic;
 signal LOCK_zd : std_ulogic;
 signal SDO_zd : std_ulogic;
 signal Violation : std_ulogic;

 -- Functional signals 
 signal not_resetb  		 : std_logic; 
 signal SPLLOUT1net, SPLLOUT2net : std_logic; 
 signal PLLOUTCOREA_temp 	 : std_logic; 
 signal PLLOUTGLOBALA_temp 	 : std_logic; 
 signal PLLOUTCOREB_temp 	 : std_logic; 
 signal PLLOUTGLOBALB_temp 	 : std_logic; 


begin 

 WireDelay   : block
 begin
          VitalWireDelay (PACKAGEPIN_ipd, PACKAGEPIN, tipd_PACKAGEPIN);
          VitalWireDelay (EXTFEEDBACK_ipd,  EXTFEEDBACK, tipd_EXTFEEDBACK);
	  DYNAMIC_DELAY : for i in 7 downto 0 generate 
	          VitalWireDelay (DYNAMICDELAY_ipd(i),DYNAMICDELAY(i),tipd_DYNAMICDELAY(i));
	  end generate DYNAMIC_DELAY; 
          VitalWireDelay (BYPASS_ipd,BYPASS, tipd_BYPASS);
          VitalWireDelay (RESETB_ipd,RESETB, tipd_RESETB);
          VitalWireDelay (SDI_ipd, SDI, tipd_SDI);
          VitalWireDelay (SCLK_ipd, SCLK, tipd_SCLK);
          VitalWireDelay (LATCHINPUTVALUE_ipd, LATCHINPUTVALUE, tipd_LATCHINPUTVALUE);
 end block;

 ------ Behavioral Section   
 not_resetb <= not(RESETB_ipd);  
 
 D: if(TEST_MODE='1') generate
 instSbtSPLL : Sbt_DS_PLL40
 generic map 	( 
		FEEDBACK_PATH 			=> FEEDBACK_PATH,
		DELAY_ADJUSTMENT_MODE_RELATIVE 	=> DELAY_ADJUSTMENT_MODE_RELATIVE,
		DELAY_ADJUSTMENT_MODE_FEEDBACK 	=> DELAY_ADJUSTMENT_MODE_FEEDBACK,
		SHIFTREG_DIV_MODE 		=> SHIFTREG_DIV_MODE,
		FDA_RELATIVE 			=> FDA_RELATIVE,
		FDA_FEEDBACK 			=> FDA_FEEDBACK,
		PLLOUT_SELECT_PORTA 		=> "GENCLK",
		PLLOUT_SELECT_PORTB 		=> PLLOUT_SELECT_PORTB, 
		DIVR 				=> DIVR,
		DIVF 				=> DIVF,
		DIVQ 				=> DIVQ,
		FILTER_RANGE 			=> FILTER_RANGE,
 		ENABLE_ICEGATE_PORTA             =>'0',
		ENABLE_ICEGATE_PORTB            =>'0' ,
        	TEST_MODE         		=> TEST_MODE
	     	)
 port map    	(
                CORE_REF_CLK 			=>open,
                EXTFEEDBACK 			=> EXTFEEDBACK_ipd,
                DYNAMICDELAY 			=> DYNAMICDELAY_ipd,
                BYPASS 				=> BYPASS_ipd,
                RESETB 				=> not_resetb ,
                PLLOUT1 			=> SPLLOUT1net,
                PLLOUT2 			=> SPLLOUT2net,
                LOCK 				=> LOCK,
                PACKAGEPIN =>PACKAGEPIN_ipd,
                PLL_SCK =>      SCLK_ipd,
                PLL_SDI =>      SDI_ipd,
                PLL_SDO =>      SDO_zd
		);
end generate D;	
 
 S: if(TEST_MODE='0') generate
instSbtSPLL : SbtSPLL40 
 generic map 	( 
		FEEDBACK_PATH 			=> FEEDBACK_PATH,
		DELAY_ADJUSTMENT_MODE_RELATIVE 	=> DELAY_ADJUSTMENT_MODE_RELATIVE,
		DELAY_ADJUSTMENT_MODE_FEEDBACK 	=> DELAY_ADJUSTMENT_MODE_FEEDBACK,
		SHIFTREG_DIV_MODE 		=> SHIFTREG_DIV_MODE,
		FDA_RELATIVE 			=> FDA_RELATIVE,
		FDA_FEEDBACK 			=> FDA_FEEDBACK,
		PLLOUT_SELECT_PORTA 		=> "GENCLK",
		PLLOUT_SELECT_PORTB 		=> PLLOUT_SELECT_PORTB, 
		DIVR 				=> DIVR,
		DIVF 				=> DIVF,
		DIVQ 				=> DIVQ,
		FILTER_RANGE 			=> FILTER_RANGE,
 		ENABLE_ICEGATE_PORTA             =>'0',
		ENABLE_ICEGATE_PORTB            =>'0' 
	     	)
 port map    	(
                REFERENCECLK 			=> PACKAGEPIN_ipd,
                EXTFEEDBACK 			=> EXTFEEDBACK_ipd,
                DYNAMICDELAY 			=> DYNAMICDELAY_ipd,
                BYPASS 				=> BYPASS_ipd,
                RESETB 				=> not_resetb ,
                PLLOUT1 			=> SPLLOUT1net,
                PLLOUT2 			=> SPLLOUT2net,
                LOCK 				=> LOCK
		);
end generate S;

  -- PLLA
 process( PLLOUTCOREA_temp, PACKAGEPIN )  
 begin 
	if(ENABLE_ICEGATE_PORTA = '1' and LATCHINPUTVALUE_ipd ='1') then 
		PLLOUTCOREA_temp <= PLLOUTCOREA_temp ; 
	else 
		PLLOUTCOREA_temp <= PACKAGEPIN; 
	end if;
 end process; 


 process( PLLOUTGLOBALA_temp, PACKAGEPIN )  
 begin 
	if(ENABLE_ICEGATE_PORTA = '1' and LATCHINPUTVALUE_ipd ='1') then 
		PLLOUTGLOBALA_temp <= PLLOUTGLOBALA_temp ; 
	else 
		PLLOUTGLOBALA_temp <= PACKAGEPIN; 
	end if; 
 end process; 

 PLLOUTCOREA_zd 	<= PLLOUTCOREA_temp; 
 PLLOUTGLOBALA_zd 	<= PLLOUTGLOBALA_temp;  

 --PLLB
 process( PLLOUTCOREB_temp, SPLLOUT2net )  
 begin 
	if(ENABLE_ICEGATE_PORTB = '1' and LATCHINPUTVALUE_ipd ='1') then 
		PLLOUTCOREB_temp <= PLLOUTCOREB_temp ; 
	else 
		PLLOUTCOREB_temp <= SPLLOUT2net; 
	end if;
 end process; 


 process( PLLOUTGLOBALB_temp, SPLLOUT2net )  
 begin 
	if(ENABLE_ICEGATE_PORTB = '1' and LATCHINPUTVALUE_ipd ='1') then 
		PLLOUTGLOBALB_temp <= PLLOUTGLOBALB_temp ; 
	else 
		PLLOUTGLOBALB_temp <= SPLLOUT2net; 
	end if; 
 end process; 

 PLLOUTCOREB_zd 	<= PLLOUTCOREB_temp; 
 PLLOUTGLOBALB_zd 	<= PLLOUTGLOBALB_temp;  
 
 VITALTimingCheck:process(SCLK_ipd,SDI_ipd)
     variable Tviol_SDI_SCLK_posedge       	: std_ulogic := '0';
     variable Tmkr_SDI_SCLK_posedge       	: VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_SDI_SCLK_negedge       	: std_ulogic := '0';
     variable Tmkr_SDI_SCLK_negedge       	: VitalTimingDataType := VitalTimingDataInit;
 begin
 if(TimingChecksOn) then
           VitalSetupHoldCheck (
        Violation      => Tviol_SDI_SCLK_posedge,
        TimingData     => Tmkr_SDI_SCLK_posedge,
        TestSignal     => SDI_ipd,
        TestSignalName => "SDI",
        TestDelay      => 0 ns,
        RefSignal      => SCLK_ipd,
        RefSignalName  => "SCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_SDI_SCLK_posedge_posedge,
        SetupLow       => tsetup_SDI_SCLK_negedge_posedge,
        HoldLow        => thold_SDI_SCLK_posedge_posedge,
        HoldHigh       => thold_SDI_SCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/PLL40",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

           VitalSetupHoldCheck (
        Violation      => Tviol_SDI_SCLK_negedge,
        TimingData     => Tmkr_SDI_SCLK_negedge,
        TestSignal     => SDI_ipd,
        TestSignalName => "SDI",
        TestDelay      => 0 ns,
        RefSignal      => SCLK_ipd,
        RefSignalName  => "SCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_SDI_SCLK_posedge_negedge,
        SetupLow       => tsetup_SDI_SCLK_negedge_negedge,
        HoldLow        => thold_SDI_SCLK_posedge_negedge,
        HoldHigh       => thold_SDI_SCLK_negedge_negedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/PLL40",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
end if;
end process VITALTimingCheck; 
 ---------------------------- 
 -- Vital Path delay  
 ---------------------------
  VITALPathDelay          : process (PLLOUTCOREA_zd, PLLOUTGLOBALA_zd,PLLOUTCOREB_zd, PLLOUTGLOBALB_zd,PACKAGEPIN_ipd,SCLK_ipd,SDO_zd )
  	variable PLLOUTCOREA_GlitchData 	: VitalGlitchDataType;
	variable PLLOUTGLOBALA_GlitchData 	: VitalGlitchDataType;
  	variable PLLOUTCOREB_GlitchData 	: VitalGlitchDataType;
	variable PLLOUTGLOBALB_GlitchData 	: VitalGlitchDataType; 
	  	variable PLLOUTCORE_GlitchData 	 : VitalGlitchDataType;
	variable PLLOUTCOREA_sig : std_ulogic := 'X';
	variable PLLOUTGLOBALA_sig : std_ulogic := 'X';	
		variable PLLOUTCOREB_sig : std_ulogic := 'X';
	variable PLLOUTGLOBALB_sig : std_ulogic := 'X';
	variable SDO_GlitchData : VitalGlitchDataType;
	variable SDO_sig : std_ulogic := 'X';
	variable LOCK_zd		 	: VitalGlitchDataType;

  begin 
	  PLLOUTCOREA_sig:=PLLOUTCOREA_zd; 
	   PLLOUTCOREB_sig:=PLLOUTCOREB_zd;
  PLLOUTGLOBALA_sig:=PLLOUTGLOBALA_zd; 
  PLLOUTGLOBALB_sig:=PLLOUTGLOBALB_zd;
  SDO_sig:=SDO_zd;
  VitalPathDelay01 (
      OutSignal                 => PLLOUTCOREA,
      GlitchData                => PLLOUTCOREA_GlitchData,
      OutSignalName             => "PLLOUTCOREA",
      OutTemp                   => PLLOUTCOREA_sig,
      Paths                     => (0 => (PACKAGEPIN_ipd'last_event, tpd_PACKAGEPIN_PLLOUTCOREA,true) ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
	  
  VitalPathDelay01 (
      OutSignal                 => PLLOUTGLOBALA,
      GlitchData                => PLLOUTGLOBALA_GlitchData,
      OutSignalName             => "PLLOUTGLOBALA",
      OutTemp                   => PLLOUTGLOBALA_sig,
      Paths                     => (0 => (PACKAGEPIN_ipd'last_event, tpd_PACKAGEPIN_PLLOUTGLOBALA, true)
									),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

  VitalPathDelay01 (
      OutSignal                 => PLLOUTCOREB,
      GlitchData                => PLLOUTCOREB_GlitchData,
      OutSignalName             => "PLLOUTCOREB",
      OutTemp                   => PLLOUTCOREB_sig,
      Paths                     => (0 => (PACKAGEPIN_ipd'last_event, tpd_PACKAGEPIN_PLLOUTCOREB,true)
							),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
	  
  VitalPathDelay01 (
      OutSignal                 => PLLOUTGLOBALB,
      GlitchData                => PLLOUTGLOBALB_GlitchData,
      OutSignalName             => "PLLOUTGLOBALB",
      OutTemp                   => PLLOUTGLOBALB_sig,
      Paths                     => (0 => (PACKAGEPIN_ipd'last_event, tpd_PACKAGEPIN_PLLOUTGLOBALB, true)
									),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
 VitalPathDelay01 (
      OutSignal                 => SDO,
      GlitchData                => SDO_GlitchData,
      OutSignalName             => "SDO",
      OutTemp                   => SDO_sig,
      Paths                     => (0 => (SCLK_ipd'last_event, tpd_SCLK_SDO_negedge, true)
									),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
  end process VITALPathDelay;	

end SB_PLL40_2_PAD_V; 


---------------------------------------------------------------------------
----			 SB_PLL40_2F_CORE 				---	
---------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;
use work.all; 

entity SB_PLL40_2F_CORE  is 
	
	generic ( 
		----------------------------------------------------------------------------------
                --VITAL PARAMETER
                ---------------------------------------------------------------------------------
                TimingChecksOn  	: boolean := true;
                Xon   			: boolean := true;
	        MsgOn 			: boolean := false;
                thold_SDI_SCLK_negedge_posedge:VitalDelayType :=0 ns;
                thold_SDI_SCLK_posedge_posedge:VitalDelayType :=0 ns;
                thold_SDI_SCLK_negedge_negedge:VitalDelayType :=0 ns;
                thold_SDI_SCLK_posedge_negedge:VitalDelayType :=0 ns;
                tsetup_SDI_SCLK_negedge_posedge:VitalDelayType :=0 ns;
                tsetup_SDI_SCLK_posedge_posedge:VitalDelayType :=0 ns;
                tsetup_SDI_SCLK_negedge_negedge:VitalDelayType :=0 ns;
                tsetup_SDI_SCLK_posedge_negedge:VitalDelayType :=0 ns; 
				tpd_SCLK_SDO_negedge          	: VitalDelayType01 := (0 ns, 0 ns);				
                --- VITAL input port delay 
                tipd_REFERENCECLK       : VitalDelayType01 := (0 ns, 0 ns);
            	tipd_EXTFEEDBACK        : VitalDelayType01 := (0 ns, 0 ns);
            	tipd_DYNAMICDELAY       : VitalDelayArrayType01(7 downto 0)  := (others => (0 ns, 0 ns));
            	tipd_BYPASS             : VitalDelayType01 := (0 ns, 0 ns);
            	tipd_RESETB             : VitalDelayType01 := (0 ns, 0 ns);
                tipd_SDI        	: VitalDelayType01 := (0 ns, 0 ns);
            	tipd_SCLK           	: VitalDelayType01 := (0 ns, 0 ns);
            	tipd_LATCHINPUTVALUE   	: VitalDelayType01 := (0 ns, 0 ns);
		-- VITAL Path Delay 	
            	tpd_REFERENCECLK_PLLOUTCOREA           	: VitalDelayType01 := (0 ns, 0 ns);
            	tpd_REFERENCECLK_PLLOUTGLOBALA          	: VitalDelayType01 := (0 ns, 0 ns);

            	tpd_REFERENCECLK_PLLOUTCOREB           	: VitalDelayType01 := (0 ns, 0 ns);
            	tpd_REFERENCECLK_PLLOUTGLOBALB          	: VitalDelayType01 := (0 ns, 0 ns);
	         -- Entity Parameters 	
		 FEEDBACK_PATH 			: string 		 :="SIMPLE";   -- SIMPLE/DELAY/PHASE_AND_DELAY/EXTERNAL 
		 DELAY_ADJUSTMENT_MODE_FEEDBACK	: string 		 :="FIXED";    -- FIXED/DYNAMIC  
		 DELAY_ADJUSTMENT_MODE_RELATIVE : string 		 :="FIXED";    -- FIXED/DYNAMIC 
		 SHIFTREG_DIV_MODE		: bit_vector(1 downto 0) := "00";      -- 00 (div by 4)/ 01 (div by 7)/11 (div by 5)   	 
		 FDA_FEEDBACK			: bit_vector(3 downto 0) :="0000";
		 FDA_RELATIVE			: bit_vector(3 downto 0) := "0000";
		 PLLOUT_SELECT_PORTA		: string 		 :="GENCLK"; 
		 PLLOUT_SELECT_PORTB		: string 		 :="GENCLK"; 

		 DIVR				: bit_vector(3 downto 0) := "0000";
		 DIVF  				: bit_vector(6 downto 0) := "0000000";
		 DIVQ	   			: bit_vector(2 downto 0) := "000";  
		 FILTER_RANGE 			: bit_vector(2 downto 0) := "000";
		 		
 		 ENABLE_ICEGATE_PORTA	        : bit 			 :='0';
 		 ENABLE_ICEGATE_PORTB	        : bit 			 :='0';
		 TEST_MODE			: bit 			 :='0';  
		 EXTERNAL_DIVIDE_FACTOR         : integer 		 := 1      -- Required for PLL Config Wizard.  
	);
	port (
                REFERENCECLK		: in std_logic;           -- PLL ref clock, driven by PAD.  
                PLLOUTCOREA	     	: out std_logic;          -- PLLA output to core logic through local routings. 
                PLLOUTGLOBALA           : out std_logic;   	  -- PLLA output to dedicated global clock network
                PLLOUTCOREB	     	: out std_logic;          -- PLLB output to core logic through local routings. 
                PLLOUTGLOBALB           : out std_logic;   	  -- PLLB output to dedicated global clock network
                EXTFEEDBACK             : in std_logic;  	  -- FB driven by core logic
                DYNAMICDELAY            : in std_logic_vector(7 downto 0);  -- driven by core logic
                LOCK                    : out std_logic;	  -- PLL Lock signal output  
                BYPASS                  : in std_logic; 	  -- REFCLK passed to PLLOUT when bypass is '1'.Driven by core logic
                RESETB                  : in std_logic; 	  -- Active low reset,Driven by core logic
                SDI                     : in std_logic;		  -- Test Input. Driven by core logic. 
                SDO                     : out std_logic; 	  -- Test output to RB Logic Tile.
                SCLK                    : in std_logic;	          -- Test Clk input.Driven by core logic. 
                LATCHINPUTVALUE         : in std_logic 		  -- iCEGate signal
	);

       attribute VITAL_LEVEL0 of SB_PLL40_2F_CORE : entity is true;

end SB_PLL40_2F_CORE; 

architecture SB_PLL40_2F_CORE_V of SB_PLL40_2F_CORE is 

	attribute VITAL_LEVEL0 of SB_PLL40_2F_CORE_V  : architecture is true;
  component Sbt_DS_PLL40  is
 
	generic ( 
		 FEEDBACK_PATH 			: string 	:="SIMPLE"; 
		 DELAY_ADJUSTMENT_MODE_FEEDBACK	: string 	:="FIXED"; 
		 DELAY_ADJUSTMENT_MODE_RELATIVE : string 	:="FIXED";
		 SHIFTREG_DIV_MODE		: bit_vector(1 downto 0) := "00"; 
		 FDA_FEEDBACK			: bit_vector(3 downto 0) :="0000";
		 FDA_RELATIVE			: bit_vector(3 downto 0) := "0000";
		 PLLOUT_SELECT_PORTA		: string 	:="GENCLK"; 
		 PLLOUT_SELECT_PORTB            : string        :="GENCLK";

		 DIVR				: bit_vector(3 downto 0) := "0000";
		 DIVF  				: bit_vector(6 downto 0) := "0000000";
		 DIVQ	   			:bit_vector(2 downto 0)  := "000";  
		 FILTER_RANGE 			:bit_vector(2 downto 0)  := "000";
		 TEST_MODE         :bit        :='0'; 		
 		ENABLE_ICEGATE_PORTA             :bit 			:='0';
		ENABLE_ICEGATE_PORTB            :bit 			:='0' 
	);
	port	(
		CORE_REF_CLK	: in    std_logic;
		EXTFEEDBACK 	: in    std_logic;
		DYNAMICDELAY	: in    std_logic_vector(7 downto 0); 
		BYPASS 		: in	std_logic;
		RESETB	 	: in 	std_logic;
		PLLOUT1 	: out  	std_logic;
		PLLOUT2		: out 	std_logic ; 
		LOCK		: out 	std_logic ;
        PACKAGEPIN : in  std_logic :='0';
        PLL_SCK     :in std_logic;
        PLL_SDI     :in std_logic;
        PLL_SDO     :out std_logic 
	); 
end component;		

 component SbtSPLL40  is
 
	generic ( 
		 FEEDBACK_PATH 			: string 	:="SIMPLE"; 
		 DELAY_ADJUSTMENT_MODE_FEEDBACK	: string 	:="FIXED"; 
		 DELAY_ADJUSTMENT_MODE_RELATIVE : string 	:="FIXED";
		 SHIFTREG_DIV_MODE		: bit_vector(1 downto 0) := "00"; 
		 FDA_FEEDBACK			: bit_vector(3 downto 0) :="0000";
		 FDA_RELATIVE			: bit_vector(3 downto 0) := "0000";
		 PLLOUT_SELECT_PORTA		: string 	:="GENCLK"; 
		 PLLOUT_SELECT_PORTB            : string        :="GENCLK"; 

		 DIVR				: bit_vector(3 downto 0) := "0000";
		 DIVF  				: bit_vector(6 downto 0) := "0000000";
		 DIVQ	   			:bit_vector(2 downto 0)  := "000";  
		 FILTER_RANGE 			:bit_vector(2 downto 0)  := "000";
		 		
 		ENABLE_ICEGATE_PORTA             :bit 			:='0';
		ENABLE_ICEGATE_PORTB            :bit 			:='0' 
	);
	port	(
		REFERENCECLK	: in    std_logic;
		EXTFEEDBACK 	: in    std_logic;
		DYNAMICDELAY	: in    std_logic_vector(7 downto 0); 
		BYPASS 		: in	std_logic;
		RESETB	 	: in 	std_logic;
		PLLOUT1 	: out  	std_logic;
		PLLOUT2		: out 	std_logic ; 
		LOCK		: out 	std_logic  
	); 
end component;

  -- Vital Wire Delay Signals   	
  signal REFERENCECLK_ipd 	: std_ulogic := 'X';
  signal EXTFEEDBACK_ipd  	: std_ulogic := 'X';
  signal DYNAMICDELAY_ipd  	: std_logic_vector(7 downto 0) := (others =>'X');
  signal BYPASS_ipd   		: std_ulogic := 'X';
  signal RESETB_ipd 		: std_ulogic := 'X';
  signal SDI_ipd  		: std_ulogic := 'X';
  signal SCLK_ipd  		: std_ulogic := 'X';
  signal LATCHINPUTVALUE_ipd  	: std_ulogic := 'X';

 -- Vital output logic signals
 signal PLLOUTCOREA_zd : std_ulogic;
 signal PLLOUTGLOBALA_zd : std_ulogic;
 signal PLLOUTCOREB_zd : std_ulogic;
 signal PLLOUTGLOBALB_zd : std_ulogic;
 signal LOCK_zd : std_ulogic;
 signal SDO_zd : std_ulogic;
 signal Violation : std_ulogic;

 -- Functional signals 
 signal not_resetb  		 : std_logic; 
 signal SPLLOUT1net, SPLLOUT2net : std_logic; 
 signal PLLOUTCOREA_temp 	 : std_logic; 
 signal PLLOUTGLOBALA_temp 	 : std_logic; 
 signal PLLOUTCOREB_temp 	 : std_logic; 
 signal PLLOUTGLOBALB_temp 	 : std_logic; 


begin 

 WireDelay   : block
 begin
          VitalWireDelay (REFERENCECLK_ipd, REFERENCECLK, tipd_REFERENCECLK);
          VitalWireDelay (EXTFEEDBACK_ipd,  EXTFEEDBACK, tipd_EXTFEEDBACK);
	  DYNAMIC_DELAY : for i in 7 downto 0 generate 
	          VitalWireDelay (DYNAMICDELAY_ipd(i),DYNAMICDELAY(i),tipd_DYNAMICDELAY(i));
	  end generate DYNAMIC_DELAY; 
          VitalWireDelay (BYPASS_ipd,BYPASS, tipd_BYPASS);
          VitalWireDelay (RESETB_ipd,RESETB, tipd_RESETB);
          VitalWireDelay (SDI_ipd, SDI, tipd_SDI);
          VitalWireDelay (SCLK_ipd, SCLK, tipd_SCLK);
          VitalWireDelay (LATCHINPUTVALUE_ipd, LATCHINPUTVALUE, tipd_LATCHINPUTVALUE);
 end block;

 ------ Behavioral Section   
 not_resetb <= not(RESETB_ipd);  
 D: if(TEST_MODE='1') generate
 instSbtSPLL : Sbt_DS_PLL40
 generic map 	( 
		FEEDBACK_PATH 			=> FEEDBACK_PATH,
		DELAY_ADJUSTMENT_MODE_RELATIVE 	=> DELAY_ADJUSTMENT_MODE_RELATIVE,
		DELAY_ADJUSTMENT_MODE_FEEDBACK 	=> DELAY_ADJUSTMENT_MODE_FEEDBACK,
		SHIFTREG_DIV_MODE 		=> SHIFTREG_DIV_MODE,
		FDA_RELATIVE 			=> FDA_RELATIVE,
		FDA_FEEDBACK 			=> FDA_FEEDBACK,
		PLLOUT_SELECT_PORTA 		=> PLLOUT_SELECT_PORTA,
		PLLOUT_SELECT_PORTB 		=> PLLOUT_SELECT_PORTB, 
		DIVR 				=> DIVR,
		DIVF 				=> DIVF,
		DIVQ 				=> DIVQ,
		FILTER_RANGE 			=> FILTER_RANGE,
 		ENABLE_ICEGATE_PORTA             =>'0',
		ENABLE_ICEGATE_PORTB            =>'0', 
        TEST_MODE          => TEST_MODE 
	     	)
 port map    	(
                CORE_REF_CLK 			=> REFERENCECLK_ipd,
                EXTFEEDBACK 			=> EXTFEEDBACK_ipd,
                DYNAMICDELAY 			=> DYNAMICDELAY_ipd,
                BYPASS 				=> BYPASS_ipd,
                RESETB 				=> not_resetb ,
                PLLOUT1 			=> SPLLOUT1net,
                PLLOUT2 			=> SPLLOUT2net,
                LOCK 				=> LOCK,
                PACKAGEPIN =>open,
                PLL_SCK =>      SCLK_ipd,
                PLL_SDI =>      SDI_ipd,
                PLL_SDO =>      SDO_zd
		);

end generate D;	  
S: if(TEST_MODE='0') generate
 instSbtSPLL : SbtSPLL40 
 generic map 	( 
		FEEDBACK_PATH 			=> FEEDBACK_PATH,
		DELAY_ADJUSTMENT_MODE_RELATIVE 	=> DELAY_ADJUSTMENT_MODE_RELATIVE,
		DELAY_ADJUSTMENT_MODE_FEEDBACK 	=> DELAY_ADJUSTMENT_MODE_FEEDBACK,
		SHIFTREG_DIV_MODE 		=> SHIFTREG_DIV_MODE,
		FDA_RELATIVE 			=> FDA_RELATIVE,
		FDA_FEEDBACK 			=> FDA_FEEDBACK,
		PLLOUT_SELECT_PORTA 		=> PLLOUT_SELECT_PORTA,
		PLLOUT_SELECT_PORTB 		=> PLLOUT_SELECT_PORTB, 
		DIVR 				=> DIVR,
		DIVF 				=> DIVF,
		DIVQ 				=> DIVQ,
		FILTER_RANGE 			=> FILTER_RANGE,
 		ENABLE_ICEGATE_PORTA             =>'0',
		ENABLE_ICEGATE_PORTB            =>'0' 
	     	)
 port map    	(
                REFERENCECLK 			=> REFERENCECLK_ipd,
                EXTFEEDBACK 			=> EXTFEEDBACK_ipd,
                DYNAMICDELAY 			=> DYNAMICDELAY_ipd,
                BYPASS 				=> BYPASS_ipd,
                RESETB 				=> not_resetb ,
                PLLOUT1 			=> SPLLOUT1net,
                PLLOUT2 			=> SPLLOUT2net,
                LOCK 				=> LOCK
		);

end generate S;	 
  -- PLLA
 process(PLLOUTCOREA_temp, SPLLOUT1net)  
 begin 
	if(ENABLE_ICEGATE_PORTA = '1' and LATCHINPUTVALUE_ipd ='1') then 
		PLLOUTCOREA_temp <= PLLOUTCOREA_temp ; 
	else 
		PLLOUTCOREA_temp <= SPLLOUT1net; 
	end if;
 end process; 


 process(PLLOUTGLOBALA_temp, SPLLOUT1net)  
 begin 
	if(ENABLE_ICEGATE_PORTA = '1' and LATCHINPUTVALUE_ipd ='1') then 
		PLLOUTGLOBALA_temp <= PLLOUTGLOBALA_temp ; 
	else 
		PLLOUTGLOBALA_temp <= SPLLOUT1net; 
	end if; 
 end process; 

 PLLOUTCOREA_zd 	<= PLLOUTCOREA_temp; 
 PLLOUTGLOBALA_zd 	<= PLLOUTGLOBALA_temp;  

 --PLLB

 process(PLLOUTCOREB_temp, SPLLOUT2net)  
 begin 
	if(ENABLE_ICEGATE_PORTB = '1' and LATCHINPUTVALUE_ipd ='1') then 
		PLLOUTCOREB_temp <= PLLOUTCOREB_temp ; 
	else 
		PLLOUTCOREB_temp <= SPLLOUT2net; 
	end if;
 end process; 


 process(PLLOUTGLOBALB_temp, SPLLOUT2net)  
 begin 
	if(ENABLE_ICEGATE_PORTB = '1' and LATCHINPUTVALUE_ipd ='1') then 
		PLLOUTGLOBALB_temp <= PLLOUTGLOBALB_temp ; 
	else 
		PLLOUTGLOBALB_temp <= SPLLOUT2net; 
	end if; 
 end process; 

 PLLOUTCOREB_zd 	<= PLLOUTCOREB_temp; 
 PLLOUTGLOBALB_zd 	<= PLLOUTGLOBALB_temp;  
 
 VITALTimingCheck:process(SCLK_ipd,SDI_ipd)
     variable Tviol_SDI_SCLK_posedge       	: std_ulogic := '0';
     variable Tmkr_SDI_SCLK_posedge       	: VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_SDI_SCLK_negedge       	: std_ulogic := '0';
     variable Tmkr_SDI_SCLK_negedge       	: VitalTimingDataType := VitalTimingDataInit;
 begin
 if(TimingChecksOn) then
           VitalSetupHoldCheck (
        Violation      => Tviol_SDI_SCLK_posedge,
        TimingData     => Tmkr_SDI_SCLK_posedge,
        TestSignal     => SDI_ipd,
        TestSignalName => "SDI",
        TestDelay      => 0 ns,
        RefSignal      => SCLK_ipd,
        RefSignalName  => "SCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_SDI_SCLK_posedge_posedge,
        SetupLow       => tsetup_SDI_SCLK_negedge_posedge,
        HoldLow        => thold_SDI_SCLK_posedge_posedge,
        HoldHigh       => thold_SDI_SCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/PLL40",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

           VitalSetupHoldCheck (
        Violation      => Tviol_SDI_SCLK_negedge,
        TimingData     => Tmkr_SDI_SCLK_negedge,
        TestSignal     => SDI_ipd,
        TestSignalName => "SDI",
        TestDelay      => 0 ns,
        RefSignal      => SCLK_ipd,
        RefSignalName  => "SCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_SDI_SCLK_posedge_negedge,
        SetupLow       => tsetup_SDI_SCLK_negedge_negedge,
        HoldLow        => thold_SDI_SCLK_posedge_negedge,
        HoldHigh       => thold_SDI_SCLK_negedge_negedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/PLL40",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
end if;
end process VITALTimingCheck; 
 ---------------------------- 
 -- Vital Path delay  
 ---------------------------
 VITALPathDelay          : process (PLLOUTCOREA_zd, PLLOUTGLOBALA_zd,PLLOUTCOREB_zd, PLLOUTGLOBALB_zd,REFERENCECLK_ipd,SCLK_ipd,SDO_zd ) 
   	variable PLLOUTCORE_GlitchData 	 : VitalGlitchDataType;
	variable PLLOUTCORE_sig : std_ulogic := 'X';
	variable PLLOUTGLOBAL_GlitchData : VitalGlitchDataType;
	variable PLLOUTGLOBAL_sig : std_ulogic := 'X';
	variable SDO_GlitchData : VitalGlitchDataType;
	variable SDO_sig : std_ulogic := 'X';
  	variable PLLOUTCOREA_GlitchData 	: VitalGlitchDataType;
	variable PLLOUTGLOBALA_GlitchData 	: VitalGlitchDataType;
  	variable PLLOUTCOREB_GlitchData 	: VitalGlitchDataType;
	variable PLLOUTGLOBALB_GlitchData 	: VitalGlitchDataType;
	variable LOCK_zd		 	: VitalGlitchDataType;
		variable PLLOUTCOREA_sig : std_ulogic := 'X';  
		variable PLLOUTCOREB_sig : std_ulogic := 'X';
	variable PLLOUTGLOBALA_sig : std_ulogic := 'X';
		variable PLLOUTGLOBALB_sig : std_ulogic := 'X';
  begin 
	  	  PLLOUTCOREA_sig:=PLLOUTCOREA_zd; 
	   PLLOUTCOREB_sig:=PLLOUTCOREB_zd;
  PLLOUTGLOBALA_sig:=PLLOUTGLOBALA_zd; 
  PLLOUTGLOBALB_sig:=PLLOUTGLOBALB_zd;
  SDO_sig:=SDO_zd;
  VitalPathDelay01 (
      OutSignal                 => PLLOUTCOREA,
      GlitchData                => PLLOUTCOREA_GlitchData,
      OutSignalName             => "PLLOUTCOREA",
      OutTemp                   => PLLOUTCOREA_zd,
      Paths                     => (0 => (REFERENCECLK_ipd'last_event, tpd_REFERENCECLK_PLLOUTCOREA,true)
							),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
	  
  VitalPathDelay01 (
      OutSignal                 => PLLOUTGLOBALA,
      GlitchData                => PLLOUTGLOBALA_GlitchData,
      OutSignalName             => "PLLOUTGLOBALA",
      OutTemp                   => PLLOUTGLOBALA_zd,
      Paths                     => (0 => (REFERENCECLK_ipd'last_event, tpd_REFERENCECLK_PLLOUTGLOBALA, true)
									),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

  VitalPathDelay01 (
      OutSignal                 => PLLOUTCOREB,
      GlitchData                => PLLOUTCOREB_GlitchData,
      OutSignalName             => "PLLOUTCOREB",
      OutTemp                   => PLLOUTCOREB_zd,
      Paths                     => (0 => (REFERENCECLK_ipd'last_event, tpd_REFERENCECLK_PLLOUTCOREB,true)
							),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
	  
  VitalPathDelay01 (
      OutSignal                 => PLLOUTGLOBALB,
      GlitchData                => PLLOUTGLOBALB_GlitchData,
      OutSignalName             => "PLLOUTGLOBALB",
      OutTemp                   => PLLOUTGLOBALB_zd,
      Paths                     => (0 => (REFERENCECLK_ipd'last_event, tpd_REFERENCECLK_PLLOUTGLOBALB, true)
									),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);  
	        VitalPathDelay01 (
      OutSignal                 => SDO,
      GlitchData                => SDO_GlitchData,
      OutSignalName             => "SDO",
      OutTemp                   => SDO_sig,
      Paths                     => (0 => (SCLK_ipd'last_event, tpd_SCLK_SDO_negedge, true)
									),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);	  
 end process VITALPathDelay;	

end SB_PLL40_2F_CORE_V;



---------------------------------------------------------------------------
----			 SB_PLL40_2F_PAD 				---	
---------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;
use work.all; 

entity SB_PLL40_2F_PAD  is 
	
	generic ( 
		----------------------------------------------------------------------------------
                --VITAL PARAMETER
                ---------------------------------------------------------------------------------
                TimingChecksOn  	: boolean := true;
                Xon   			: boolean := true;
	        MsgOn 			: boolean := false;	
                thold_SDI_SCLK_negedge_posedge:VitalDelayType :=0 ns;
                thold_SDI_SCLK_posedge_posedge:VitalDelayType :=0 ns;
                thold_SDI_SCLK_negedge_negedge:VitalDelayType :=0 ns;
                thold_SDI_SCLK_posedge_negedge:VitalDelayType :=0 ns;
                tsetup_SDI_SCLK_negedge_posedge:VitalDelayType :=0 ns;
                tsetup_SDI_SCLK_posedge_posedge:VitalDelayType :=0 ns;
                tsetup_SDI_SCLK_negedge_negedge:VitalDelayType :=0 ns;
                tsetup_SDI_SCLK_posedge_negedge:VitalDelayType :=0 ns; 
				tpd_SCLK_SDO_negedge          	: VitalDelayType01 := (0 ns, 0 ns);	
                --- VITAL input port delay 
                tipd_PACKAGEPIN       : VitalDelayType01 := (0 ns, 0 ns);
            	tipd_EXTFEEDBACK        : VitalDelayType01 := (0 ns, 0 ns);
            	tipd_DYNAMICDELAY       : VitalDelayArrayType01(7 downto 0)  := (others => (0 ns, 0 ns));
            	tipd_BYPASS             : VitalDelayType01 := (0 ns, 0 ns);
            	tipd_RESETB             : VitalDelayType01 := (0 ns, 0 ns);
                tipd_SDI        	: VitalDelayType01 := (0 ns, 0 ns);
            	tipd_SCLK           	: VitalDelayType01 := (0 ns, 0 ns);
            	tipd_LATCHINPUTVALUE   	: VitalDelayType01 := (0 ns, 0 ns);
		-- VITAL Path Delay 	
            	tpd_PACKAGEPIN_PLLOUTCOREA           	: VitalDelayType01 := (0 ns, 0 ns);
            	tpd_PACKAGEPIN_PLLOUTGLOBALA          	: VitalDelayType01 := (0 ns, 0 ns);

            	tpd_PACKAGEPIN_PLLOUTCOREB           	: VitalDelayType01 := (0 ns, 0 ns);
            	tpd_PACKAGEPIN_PLLOUTGLOBALB          	: VitalDelayType01 := (0 ns, 0 ns);
	         -- Entity Parameters 	
		 FEEDBACK_PATH 			: string 		 :="SIMPLE";   -- SIMPLE/DELAY/PHASE_AND_DELAY/EXTERNAL 
		 DELAY_ADJUSTMENT_MODE_FEEDBACK	: string 		 :="FIXED";    -- FIXED/DYNAMIC  
		 DELAY_ADJUSTMENT_MODE_RELATIVE : string 		 :="FIXED";    -- FIXED/DYNAMIC 
		 SHIFTREG_DIV_MODE		:  bit_vector(1 downto 0) := "00";      -- 00 (div by 4)/ 01 (div by 7)/11 (div by 5)   	 
		 FDA_FEEDBACK			: bit_vector(3 downto 0) :="0000";
		 FDA_RELATIVE			: bit_vector(3 downto 0) := "0000";
		 PLLOUT_SELECT_PORTA		: string 		 :="GENCLK"; 
		 PLLOUT_SELECT_PORTB		: string 		 :="GENCLK"; 

		 DIVR				: bit_vector(3 downto 0) := "0000";
		 DIVF  				: bit_vector(6 downto 0) := "0000000";
		 DIVQ	   			: bit_vector(2 downto 0) := "000";  
		 FILTER_RANGE 			: bit_vector(2 downto 0) := "000";
		 		
 		 ENABLE_ICEGATE_PORTA	        : bit 			 :='0';
 		 ENABLE_ICEGATE_PORTB	        : bit 			 :='0';
		 TEST_MODE			: bit 			 :='0';  
		 EXTERNAL_DIVIDE_FACTOR         : integer 		 := 1      -- Required for PLL Config Wizard.  
	);
	port (
                PACKAGEPIN		: in std_logic;           -- PLL ref clock, driven by PAD.  
                PLLOUTCOREA	     	: out std_logic;          -- PLLA output to core logic through local routings. 
                PLLOUTGLOBALA           : out std_logic;   	  -- PLLA output to dedicated global clock network
                PLLOUTCOREB	     	: out std_logic;          -- PLLB output to core logic through local routings. 
                PLLOUTGLOBALB           : out std_logic;   	  -- PLLB output to dedicated global clock network
                EXTFEEDBACK             : in std_logic;  	  -- FB driven by core logic
                DYNAMICDELAY            : in std_logic_vector(7 downto 0);  -- driven by core logic
                LOCK                    : out std_logic;	  -- PLL Lock signal output  
                BYPASS                  : in std_logic; 	  -- REFCLK passed to PLLOUT when bypass is '1'.Driven by core logic
                RESETB                  : in std_logic; 	  -- Active low reset,Driven by core logic
                SDI                     : in std_logic;		  -- Test Input. Driven by core logic. 
                SDO                     : out std_logic; 	  -- Test output to RB Logic Tile.
                SCLK                    : in std_logic;	          -- Test Clk input.Driven by core logic. 
                LATCHINPUTVALUE         : in std_logic 		  -- iCEGate signal
	);

       attribute VITAL_LEVEL0 of SB_PLL40_2F_PAD : entity is true;

end SB_PLL40_2F_PAD; 

architecture SB_PLL40_2F_PAD_V of SB_PLL40_2F_PAD is 

	attribute VITAL_LEVEL0 of SB_PLL40_2F_PAD_V  : architecture is true;
 component Sbt_DS_PLL40  is
 
	generic ( 
		 FEEDBACK_PATH 			: string 	:="SIMPLE"; 
		 DELAY_ADJUSTMENT_MODE_FEEDBACK	: string 	:="FIXED"; 
		 DELAY_ADJUSTMENT_MODE_RELATIVE : string 	:="FIXED";
		 SHIFTREG_DIV_MODE		: bit_vector(1 downto 0) := "00"; 
		 FDA_FEEDBACK			: bit_vector(3 downto 0) :="0000";
		 FDA_RELATIVE			: bit_vector(3 downto 0) := "0000";
		 PLLOUT_SELECT_PORTA		: string 	:="GENCLK"; 
		 PLLOUT_SELECT_PORTB            : string        :="GENCLK";

		 DIVR				: bit_vector(3 downto 0) := "0000";
		 DIVF  				: bit_vector(6 downto 0) := "0000000";
		 DIVQ	   			:bit_vector(2 downto 0)  := "000";  
		 FILTER_RANGE 			:bit_vector(2 downto 0)  := "000";
		 TEST_MODE         :bit        :='0'; 		
 		ENABLE_ICEGATE_PORTA             :bit 			:='0';
		ENABLE_ICEGATE_PORTB            :bit 			:='0' 
	);
	port	(
		CORE_REF_CLK	: in    std_logic:='0';
		EXTFEEDBACK 	: in    std_logic;
		DYNAMICDELAY	: in    std_logic_vector(7 downto 0); 
		BYPASS 		: in	std_logic;
		RESETB	 	: in 	std_logic;
		PLLOUT1 	: out  	std_logic;
		PLLOUT2		: out 	std_logic ; 
		LOCK		: out 	std_logic ;
        PACKAGEPIN : in  std_logic :='0';
        PLL_SCK     :in std_logic;
        PLL_SDI     :in std_logic;
        PLL_SDO     :out std_logic 
	); 
end component;	

 component SbtSPLL40  is
 
	generic ( 
		 FEEDBACK_PATH 			: string 	:="SIMPLE"; 
		 DELAY_ADJUSTMENT_MODE_FEEDBACK	: string 	:="FIXED"; 
		 DELAY_ADJUSTMENT_MODE_RELATIVE : string 	:="FIXED";
		 SHIFTREG_DIV_MODE		: bit_vector(1 downto 0) := "00"; 
		 FDA_FEEDBACK			: bit_vector(3 downto 0) :="0000";
		 FDA_RELATIVE			: bit_vector(3 downto 0) := "0000";
		 PLLOUT_SELECT_PORTA		: string 	:="GENCLK"; 
		 PLLOUT_SELECT_PORTB            : string        :="GENCLK"; 

		 DIVR				: bit_vector(3 downto 0) := "0000";
		 DIVF  				: bit_vector(6 downto 0) := "0000000";
		 DIVQ	   			:bit_vector(2 downto 0)  := "000";  
		 FILTER_RANGE 			:bit_vector(2 downto 0)  := "000";
		 		
 		ENABLE_ICEGATE_PORTA             :bit 			:='0';
		ENABLE_ICEGATE_PORTB            :bit 			:='0' 
	);
	port	(
		REFERENCECLK	: in    std_logic;
		EXTFEEDBACK 	: in    std_logic;
		DYNAMICDELAY	: in    std_logic_vector(7 downto 0); 
		BYPASS 		: in	std_logic;
		RESETB	 	: in 	std_logic;
		PLLOUT1 	: out  	std_logic;
		PLLOUT2		: out 	std_logic ; 
		LOCK		: out 	std_logic  
	); 
end component;

  -- Vital Wire Delay Signals   	
  signal PACKAGEPIN_ipd 	: std_ulogic := 'X';
  signal EXTFEEDBACK_ipd  	: std_ulogic := 'X';
  signal DYNAMICDELAY_ipd  	: std_logic_vector(7 downto 0) := (others =>'X');
  signal BYPASS_ipd   		: std_ulogic := 'X';
  signal RESETB_ipd 		: std_ulogic := 'X';
  signal SDI_ipd  		: std_ulogic := 'X';
  signal SCLK_ipd  		: std_ulogic := 'X';
  signal LATCHINPUTVALUE_ipd  	: std_ulogic := 'X';

 -- Vital output logic signals
 signal PLLOUTCOREA_zd : std_ulogic;
 signal PLLOUTGLOBALA_zd : std_ulogic;
 signal PLLOUTCOREB_zd : std_ulogic;
 signal PLLOUTGLOBALB_zd : std_ulogic;
 signal LOCK_zd : std_ulogic;
 signal SDO_zd : std_ulogic;
 signal Violation : std_ulogic;

 -- Functional signals 
 signal not_resetb  		 : std_logic; 
 signal SPLLOUT1net, SPLLOUT2net : std_logic; 
 signal PLLOUTCOREA_temp 	 : std_logic; 
 signal PLLOUTGLOBALA_temp 	 : std_logic; 
 signal PLLOUTCOREB_temp 	 : std_logic; 
 signal PLLOUTGLOBALB_temp 	 : std_logic; 


begin 

 WireDelay   : block
 begin
          VitalWireDelay (PACKAGEPIN_ipd, PACKAGEPIN, tipd_PACKAGEPIN);
          VitalWireDelay (EXTFEEDBACK_ipd,  EXTFEEDBACK, tipd_EXTFEEDBACK);
	  DYNAMIC_DELAY : for i in 7 downto 0 generate 
	          VitalWireDelay (DYNAMICDELAY_ipd(i),DYNAMICDELAY(i),tipd_DYNAMICDELAY(i));
	  end generate DYNAMIC_DELAY; 
          VitalWireDelay (BYPASS_ipd,BYPASS, tipd_BYPASS);
          VitalWireDelay (RESETB_ipd,RESETB, tipd_RESETB);
          VitalWireDelay (SDI_ipd, SDI, tipd_SDI);
          VitalWireDelay (SCLK_ipd, SCLK, tipd_SCLK);
          VitalWireDelay (LATCHINPUTVALUE_ipd, LATCHINPUTVALUE, tipd_LATCHINPUTVALUE);
 end block;

 ------ Behavioral Section   
 not_resetb <= not(RESETB_ipd);  
 
 D: if(TEST_MODE='1') generate
 instSbtSPLL : Sbt_DS_PLL40
 generic map 	( 
		FEEDBACK_PATH 			=> FEEDBACK_PATH,
		DELAY_ADJUSTMENT_MODE_RELATIVE 	=> DELAY_ADJUSTMENT_MODE_RELATIVE,
		DELAY_ADJUSTMENT_MODE_FEEDBACK 	=> DELAY_ADJUSTMENT_MODE_FEEDBACK,
		SHIFTREG_DIV_MODE 		=> SHIFTREG_DIV_MODE,
		FDA_RELATIVE 			=> FDA_RELATIVE,
		FDA_FEEDBACK 			=> FDA_FEEDBACK,
		PLLOUT_SELECT_PORTA 		=> PLLOUT_SELECT_PORTA,
		PLLOUT_SELECT_PORTB 		=> PLLOUT_SELECT_PORTB, 
		DIVR 				=> DIVR,
		DIVF 				=> DIVF,
		DIVQ 				=> DIVQ,
		FILTER_RANGE 			=> FILTER_RANGE,
 		ENABLE_ICEGATE_PORTA             =>'0',
		ENABLE_ICEGATE_PORTB            =>'0' ,
        TEST_MODE          => TEST_MODE
	     	)
 port map    	(
                CORE_REF_CLK 			=>open,
                EXTFEEDBACK 			=> EXTFEEDBACK_ipd,
                DYNAMICDELAY 			=> DYNAMICDELAY_ipd,
                BYPASS 				=> BYPASS_ipd,
                RESETB 				=> not_resetb ,
                PLLOUT1 			=> SPLLOUT1net,
                PLLOUT2 			=> SPLLOUT2net,
                LOCK 				=> LOCK,
                PACKAGEPIN =>PACKAGEPIN_ipd,
                PLL_SCK =>      SCLK_ipd,
                PLL_SDI =>      SDI_ipd,
                PLL_SDO =>      SDO_zd
		);
end generate D;	
 
S: if(TEST_MODE='0') generate
instSbtSPLL : SbtSPLL40 
 generic map 	( 
		FEEDBACK_PATH 			=> FEEDBACK_PATH,
		DELAY_ADJUSTMENT_MODE_RELATIVE 	=> DELAY_ADJUSTMENT_MODE_RELATIVE,
		DELAY_ADJUSTMENT_MODE_FEEDBACK 	=> DELAY_ADJUSTMENT_MODE_FEEDBACK,
		SHIFTREG_DIV_MODE 		=> SHIFTREG_DIV_MODE,
		FDA_RELATIVE 			=> FDA_RELATIVE,
		FDA_FEEDBACK 			=> FDA_FEEDBACK,
		PLLOUT_SELECT_PORTA 		=> PLLOUT_SELECT_PORTA,
		PLLOUT_SELECT_PORTB 		=> PLLOUT_SELECT_PORTB, 
		DIVR 				=> DIVR,
		DIVF 				=> DIVF,
		DIVQ 				=> DIVQ,
		FILTER_RANGE 			=> FILTER_RANGE,
 		ENABLE_ICEGATE_PORTA             =>'0',
		ENABLE_ICEGATE_PORTB            =>'0' 
	     	)
 port map    	(
                REFERENCECLK 			=> PACKAGEPIN_ipd,
                EXTFEEDBACK 			=> EXTFEEDBACK_ipd,
                DYNAMICDELAY 			=> DYNAMICDELAY_ipd,
                BYPASS 				=> BYPASS_ipd,
                RESETB 				=> not_resetb ,
                PLLOUT1 			=> SPLLOUT1net,
                PLLOUT2 			=> SPLLOUT2net,
                LOCK 				=> LOCK
		);
end generate S;	

  -- PLLA
 process(PLLOUTCOREA_temp, SPLLOUT1net)  
 begin 
	if(ENABLE_ICEGATE_PORTA = '1' and LATCHINPUTVALUE_ipd ='1') then 
		PLLOUTCOREA_temp <= PLLOUTCOREA_temp ; 
	else 
		PLLOUTCOREA_temp <= SPLLOUT1net; 
	end if;
 end process; 


 process(PLLOUTGLOBALA_temp, SPLLOUT1net)  
 begin 
	if(ENABLE_ICEGATE_PORTA = '1' and LATCHINPUTVALUE_ipd ='1') then 
		PLLOUTGLOBALA_temp <= PLLOUTGLOBALA_temp ; 
	else 
		PLLOUTGLOBALA_temp <= SPLLOUT1net; 
	end if; 
 end process; 

 PLLOUTCOREA_zd 	<= PLLOUTCOREA_temp; 
 PLLOUTGLOBALA_zd 	<= PLLOUTGLOBALA_temp;  

 --PLLB

 process(PLLOUTCOREB_temp, SPLLOUT2net)  
 begin 
	if(ENABLE_ICEGATE_PORTB = '1' and LATCHINPUTVALUE_ipd ='1') then 
		PLLOUTCOREB_temp <= PLLOUTCOREB_temp ; 
	else 
		PLLOUTCOREB_temp <= SPLLOUT2net; 
	end if;
 end process; 


 process(PLLOUTGLOBALB_temp, SPLLOUT2net)  
 begin 
	if(ENABLE_ICEGATE_PORTB = '1' and LATCHINPUTVALUE_ipd ='1') then 
		PLLOUTGLOBALB_temp <= PLLOUTGLOBALB_temp ; 
	else 
		PLLOUTGLOBALB_temp <= SPLLOUT2net; 
	end if; 
 end process; 

 PLLOUTCOREB_zd 	<= PLLOUTCOREB_temp; 
 PLLOUTGLOBALB_zd 	<= PLLOUTGLOBALB_temp;  

  VITALTimingCheck:process(SCLK_ipd,SDI_ipd)
     variable Tviol_SDI_SCLK_posedge       	: std_ulogic := '0';
     variable Tmkr_SDI_SCLK_posedge       	: VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_SDI_SCLK_negedge       	: std_ulogic := '0';
     variable Tmkr_SDI_SCLK_negedge       	: VitalTimingDataType := VitalTimingDataInit;
 begin
 if(TimingChecksOn) then
           VitalSetupHoldCheck (
        Violation      => Tviol_SDI_SCLK_posedge,
        TimingData     => Tmkr_SDI_SCLK_posedge,
        TestSignal     => SDI_ipd,
        TestSignalName => "SDI",
        TestDelay      => 0 ns,
        RefSignal      => SCLK_ipd,
        RefSignalName  => "SCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_SDI_SCLK_posedge_posedge,
        SetupLow       => tsetup_SDI_SCLK_negedge_posedge,
        HoldLow        => thold_SDI_SCLK_posedge_posedge,
        HoldHigh       => thold_SDI_SCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/PLL40",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

           VitalSetupHoldCheck (
        Violation      => Tviol_SDI_SCLK_negedge,
        TimingData     => Tmkr_SDI_SCLK_negedge,
        TestSignal     => SDI_ipd,
        TestSignalName => "SDI",
        TestDelay      => 0 ns,
        RefSignal      => SCLK_ipd,
        RefSignalName  => "SCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_SDI_SCLK_posedge_negedge,
        SetupLow       => tsetup_SDI_SCLK_negedge_negedge,
        HoldLow        => thold_SDI_SCLK_posedge_negedge,
        HoldHigh       => thold_SDI_SCLK_negedge_negedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/PLL40",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
end if;
end process VITALTimingCheck;
 ---------------------------- 
 -- Vital Path delay  
 ---------------------------
 VITALPathDelay          : process (PLLOUTCOREA_zd, PLLOUTGLOBALA_zd,PLLOUTCOREB_zd, PLLOUTGLOBALB_zd,PACKAGEPIN_ipd,SCLK_ipd,SDO_zd)	   
   	variable PLLOUTCORE_GlitchData 	 : VitalGlitchDataType;
	variable PLLOUTCOREA_sig : std_ulogic := 'X';  
		variable PLLOUTCOREB_sig : std_ulogic := 'X';
	variable PLLOUTGLOBALA_sig : std_ulogic := 'X';
		variable PLLOUTGLOBALB_sig : std_ulogic := 'X';
	variable SDO_GlitchData : VitalGlitchDataType;
	variable SDO_sig : std_ulogic := 'X';
  	variable PLLOUTCOREA_GlitchData 	: VitalGlitchDataType;
	variable PLLOUTGLOBALA_GlitchData 	: VitalGlitchDataType;
  	variable PLLOUTCOREB_GlitchData 	: VitalGlitchDataType;
	variable PLLOUTGLOBALB_GlitchData 	: VitalGlitchDataType;
	variable LOCK_zd		 	: VitalGlitchDataType;

  begin
	  PLLOUTCOREA_sig:=PLLOUTCOREA_zd; 
	   PLLOUTCOREB_sig:=PLLOUTCOREB_zd;
  PLLOUTGLOBALA_sig:=PLLOUTGLOBALA_zd; 
  PLLOUTGLOBALB_sig:=PLLOUTGLOBALB_zd;
  SDO_sig:=SDO_zd;
  VitalPathDelay01 (
      OutSignal                 => PLLOUTCOREA,
      GlitchData                => PLLOUTCOREA_GlitchData,
      OutSignalName             => "PLLOUTCOREA",
      OutTemp                   => PLLOUTCOREA_sig,
      Paths                     => (0 => (PACKAGEPIN_ipd'last_event, tpd_PACKAGEPIN_PLLOUTCOREA,true)
							),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
	  
  VitalPathDelay01 (
      OutSignal                 => PLLOUTGLOBALA,
      GlitchData                => PLLOUTGLOBALA_GlitchData,
      OutSignalName             => "PLLOUTGLOBALA",
      OutTemp                   => PLLOUTGLOBALA_sig,
      Paths                     => (0 => (PACKAGEPIN_ipd'last_event, tpd_PACKAGEPIN_PLLOUTGLOBALA, true)
									),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

  VitalPathDelay01 (
      OutSignal                 => PLLOUTCOREB,
      GlitchData                => PLLOUTCOREB_GlitchData,
      OutSignalName             => "PLLOUTCOREB",
      OutTemp                   => PLLOUTCOREB_sig,
      Paths                     => (0 => (PACKAGEPIN_ipd'last_event, tpd_PACKAGEPIN_PLLOUTCOREB,true)
							),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
	  
  VitalPathDelay01 (
      OutSignal                 => PLLOUTGLOBALB,
      GlitchData                => PLLOUTGLOBALB_GlitchData,
      OutSignalName             => "PLLOUTGLOBALB",
      OutTemp                   => PLLOUTGLOBALB_sig,
      Paths                     => (0 => (PACKAGEPIN_ipd'last_event, tpd_PACKAGEPIN_PLLOUTGLOBALB, true)
									),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);	 
	        VitalPathDelay01 (
      OutSignal                 => SDO,
      GlitchData                => SDO_GlitchData,
      OutSignalName             => "SDO",
      OutTemp                   => SDO_sig,
      Paths                     => (0 => (SCLK_ipd'last_event, tpd_SCLK_SDO_negedge, true)
									),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
 end process VITALPathDelay;	

end SB_PLL40_2F_PAD_V; 

---------------------------------------------------------------------------
----			 SB_PLL40_PAD_DS 				---	
---------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;
use work.all; 

entity SB_PLL40_PAD_DS  is 
	
	generic ( 
		----------------------------------------------------------------------------------
                --VITAL PARAMETER
                ---------------------------------------------------------------------------------
                TimingChecksOn  	: boolean := true;
                Xon   			: boolean := true;
	        MsgOn 			: boolean := false;
                --- VITAL input port delay 
                tipd_PACKAGEPIN         : VitalDelayType01 := (0 ns, 0 ns);
                tipd_PACKAGEPINB        : VitalDelayType01 := (0 ns, 0 ns);
            	tipd_EXTFEEDBACK        : VitalDelayType01 := (0 ns, 0 ns);
            	tipd_DYNAMICDELAY       : VitalDelayArrayType01(7 downto 0)  := (others => (0 ns, 0 ns));
            	tipd_BYPASS             : VitalDelayType01 := (0 ns, 0 ns);
            	tipd_RESETB             : VitalDelayType01 := (0 ns, 0 ns);
                tipd_SDI        	: VitalDelayType01 := (0 ns, 0 ns);
            	tipd_SCLK           	: VitalDelayType01 := (0 ns, 0 ns);
            	tipd_LATCHINPUTVALUE   	: VitalDelayType01 := (0 ns, 0 ns);
		-- VITAL Path Delay 	
            	tpd_PACKAGEPIN_PLLOUTCORE           	: VitalDelayType01 := (0 ns, 0 ns);
            	tpd_PACKAGEPIN_PLLOUTGLOBAL          	: VitalDelayType01 := (0 ns, 0 ns);
	         -- Entity Parameters 	
		 FEEDBACK_PATH 			: string 		 :="SIMPLE";   -- SIMPLE/DELAY/PHASE_AND_DELAY/EXTERNAL 
		 DELAY_ADJUSTMENT_MODE_FEEDBACK	: string 		 :="FIXED";    -- FIXED/DYNAMIC  
		 DELAY_ADJUSTMENT_MODE_RELATIVE : string 		 :="FIXED";    -- FIXED/DYNAMIC 
		 SHIFTREG_DIV_MODE		:  bit_vector(1 downto 0) := "00";     -- 00 (div by 4)/ 01 (div by 7)/11 (div by 5)   	 
		 FDA_FEEDBACK			: bit_vector(3 downto 0) :="0000";
		 FDA_RELATIVE			: bit_vector(3 downto 0) := "0000";
		 PLLOUT_SELECT			: string 		 :="GENCLK"; 

		 DIVR				: bit_vector(3 downto 0) := "0000";
		 DIVF  				: bit_vector(6 downto 0) := "0000000";
		 DIVQ	   			: bit_vector(2 downto 0) := "000";  
		 FILTER_RANGE 			: bit_vector(2 downto 0) := "000";
		 		
 		 ENABLE_ICEGATE		        : bit 			 :='0';
		 TEST_MODE			: bit 			 :='0';  
		 EXTERNAL_DIVIDE_FACTOR         : integer 		 := 1      -- Required for PLL Config Wizard.  
	);
	port (
                PACKAGEPIN		: in std_logic;           -- PLL ref clock(+), driven by PAD.  
                PACKAGEPINB		: in std_logic;           -- PLL ref clock(-), driven by PAD.  
                PLLOUTCORE	     	: out std_logic;          -- PLL output to core logic through local routings. 
                PLLOUTGLOBAL            : out std_logic;   	  -- PLL output to dedicated global clock network
                EXTFEEDBACK             : in std_logic;  	  -- FB driven by core logic
                DYNAMICDELAY            : in std_logic_vector(7 downto 0);  -- driven by core logic
                LOCK                    : out std_logic;	  -- PLL Lock signal output  
                BYPASS                  : in std_logic; 	  -- REFCLK passed to PLLOUT when bypass is '1'.Driven by core logic
                RESETB                  : in std_logic; 	  -- Active low reset,Driven by core logic
                SDI                     : in std_logic;		  -- Test Input. Driven by core logic. 
                SDO                     : out std_logic; 	  -- Test output to RB Logic Tile.
                SCLK                    : in std_logic;	          -- Test Clk input.Driven by core logic. 
                LATCHINPUTVALUE         : in std_logic 		  -- iCEGate signal
	);

       attribute VITAL_LEVEL0 of SB_PLL40_PAD_DS : entity is true;

end SB_PLL40_PAD_DS; 

architecture SB_PLL40_PAD_DS_V of SB_PLL40_PAD_DS is 

	attribute VITAL_LEVEL0 of SB_PLL40_PAD_DS_V  : architecture is true;


 component SbtSPLL40  is
 
	generic ( 
		 FEEDBACK_PATH 			: string 	:="SIMPLE"; 
		 DELAY_ADJUSTMENT_MODE_FEEDBACK	: string 	:="FIXED"; 
		 DELAY_ADJUSTMENT_MODE_RELATIVE : string 	:="FIXED";
		 SHIFTREG_DIV_MODE		: bit_vector(1 downto 0) := "00"; 
		 FDA_FEEDBACK			: bit_vector(3 downto 0) :="0000";
		 FDA_RELATIVE			: bit_vector(3 downto 0) := "0000";
		 PLLOUT_SELECT_PORTA		: string 	:="GENCLK"; 
		 PLLOUT_SELECT_PORTB            : string        :="GENCLK";

		 DIVR				: bit_vector(3 downto 0) := "0000";
		 DIVF  				: bit_vector(6 downto 0) := "0000000";
		 DIVQ	   			:bit_vector(2 downto 0)  := "000";  
		 FILTER_RANGE 			:bit_vector(2 downto 0)  := "000";
		 		
 		ENABLE_ICEGATE_PORTA             :bit 			:='0';
		ENABLE_ICEGATE_PORTB            :bit 			:='0' 
	);
	port	(
		REFERENCECLK	: in    std_logic;
		EXTFEEDBACK 	: in    std_logic;
		DYNAMICDELAY	: in    std_logic_vector(7 downto 0); 
		BYPASS 		: in	std_logic;
		RESETB	 	: in 	std_logic;
		PLLOUT1 	: out  	std_logic;
		PLLOUT2		: out 	std_logic ; 
		LOCK		: out 	std_logic  
	); 
end component;

  -- Vital Wire Delay Signals   	
  signal PACKAGEPIN_ipd 	: std_ulogic := 'X';
  signal PACKAGEPINB_ipd 	: std_ulogic := 'X';
  signal EXTFEEDBACK_ipd  	: std_ulogic := 'X';
  signal DYNAMICDELAY_ipd  	: std_logic_vector(7 downto 0) := (others =>'X');
  signal BYPASS_ipd   		: std_ulogic := 'X';
  signal RESETB_ipd 		: std_ulogic := 'X';
  signal SDI_ipd  		: std_ulogic := 'X';
  signal SCLK_ipd  		: std_ulogic := 'X';
  signal LATCHINPUTVALUE_ipd  	: std_ulogic := 'X';

 -- Vital output logic signals
 signal PLLOUTCORE_zd : std_ulogic;
 signal PLLOUTGLOBAL_zd : std_ulogic;
 signal LOCK_zd : std_ulogic;
 signal SDO_zd : std_ulogic;
 signal Violation : std_ulogic;

 -- Functional Signals 
 signal not_resetb  		 : std_logic; 
 signal SPLLOUT1net, SPLLOUT2net : std_logic; 
 signal PLLOUTCORE_temp 	 : std_logic; 
 signal PLLOUTGLOBAL_temp 	 : std_logic; 

begin 

 WireDelay   : block
 begin
          VitalWireDelay (PACKAGEPIN_ipd, PACKAGEPIN, tipd_PACKAGEPIN);
          VitalWireDelay (PACKAGEPINB_ipd, PACKAGEPINB, tipd_PACKAGEPINB);
          VitalWireDelay (EXTFEEDBACK_ipd,  EXTFEEDBACK, tipd_EXTFEEDBACK);
	  DYNAMIC_DELAY : for i in 7 downto 0 generate 
	          VitalWireDelay (DYNAMICDELAY_ipd(i),DYNAMICDELAY(i),tipd_DYNAMICDELAY(i));
	  end generate DYNAMIC_DELAY; 
          VitalWireDelay (BYPASS_ipd,BYPASS, tipd_BYPASS);
          VitalWireDelay (RESETB_ipd,RESETB, tipd_RESETB);
          VitalWireDelay (SDI_ipd, SDI, tipd_SDI);
          VitalWireDelay (SCLK_ipd, SCLK, tipd_SCLK);
          VitalWireDelay (LATCHINPUTVALUE_ipd, LATCHINPUTVALUE, tipd_LATCHINPUTVALUE);
 end block;

 ------ Behavioral Section   
 not_resetb <= not(RESETB_ipd);  

 instSbtSPLL : SbtSPLL40 
 generic map 	( 
		FEEDBACK_PATH 			=> FEEDBACK_PATH,
		DELAY_ADJUSTMENT_MODE_RELATIVE 	=> DELAY_ADJUSTMENT_MODE_RELATIVE,
		DELAY_ADJUSTMENT_MODE_FEEDBACK 	=> DELAY_ADJUSTMENT_MODE_FEEDBACK,
		SHIFTREG_DIV_MODE 		=> SHIFTREG_DIV_MODE,
		FDA_RELATIVE 			=> FDA_RELATIVE,
		FDA_FEEDBACK 			=> FDA_FEEDBACK,
		PLLOUT_SELECT_PORTA 		=> PLLOUT_SELECT,
		PLLOUT_SELECT_PORTB 		=> "GENCLK",
		DIVR 				=> DIVR,
		DIVF 				=> DIVF,
		DIVQ 				=> DIVQ,
		FILTER_RANGE 			=> FILTER_RANGE,
 		ENABLE_ICEGATE_PORTA             =>'0',
		ENABLE_ICEGATE_PORTB            =>'0' 
	     	)
 port map    	(
                REFERENCECLK 			=> PACKAGEPIN_ipd,
                EXTFEEDBACK 			=> EXTFEEDBACK_ipd,
                DYNAMICDELAY 			=> DYNAMICDELAY_ipd,
                BYPASS 				=> BYPASS_ipd,
                RESETB 				=> not_resetb ,
                PLLOUT1 			=> SPLLOUT1net,
                PLLOUT2 			=> SPLLOUT2net,
                LOCK 				=> LOCK
		);



 process(PLLOUTCORE_temp, SPLLOUT1net)  
 begin 
	if(ENABLE_ICEGATE = '1' and LATCHINPUTVALUE_ipd ='1') then 
		PLLOUTCORE_temp <= PLLOUTCORE_temp ; 
	else 
		PLLOUTCORE_temp <= SPLLOUT1net; 
	end if;
 end process; 


 process(PLLOUTGLOBAL_temp, SPLLOUT1net)  
 begin 
	if(ENABLE_ICEGATE = '1' and LATCHINPUTVALUE_ipd ='1') then 
		PLLOUTGLOBAL_temp <= PLLOUTGLOBAL_temp ; 
	else 
		PLLOUTGLOBAL_temp <= SPLLOUT1net; 
	end if; 
 end process; 

 PLLOUTCORE_zd 	<= PLLOUTCORE_temp; 
 PLLOUTGLOBAL_zd 	<= PLLOUTGLOBAL_temp;  

 
 ---------------------------- 
 -- Vital Path delay  
 ---------------------------
  VITALPathDelay          : process (PLLOUTCORE_zd, PLLOUTGLOBAL_zd, PACKAGEPIN_ipd )
  	variable PLLOUTCORE_GlitchData 	 : VitalGlitchDataType;
	variable PLLOUTGLOBAL_GlitchData : VitalGlitchDataType;
	variable LOCK_zd		 : VitalGlitchDataType;

  begin 		
  VitalPathDelay01 (
      OutSignal                 => PLLOUTCORE,
      GlitchData                => PLLOUTCORE_GlitchData,
      OutSignalName             => "PLLOUTCORE",
      OutTemp                   => PLLOUTCORE_zd,
      Paths                     => (0 => (PACKAGEPIN_ipd'last_event, tpd_PACKAGEPIN_PLLOUTCORE,true)
							),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
	  
      VitalPathDelay01 (
      OutSignal                 => PLLOUTGLOBAL,
      GlitchData                => PLLOUTGLOBAL_GlitchData,
      OutSignalName             => "PLLOUTGLOBAL",
      OutTemp                   => PLLOUTGLOBAL_zd,
      Paths                     => (0 => (PACKAGEPIN_ipd'last_event, tpd_PACKAGEPIN_PLLOUTGLOBAL, true)
									),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
 end process VITALPathDelay;	

end SB_PLL40_PAD_DS_V; 


---------------------------------------------------------------------------
----			 SB_PLL40_2F_PAD_DS 				---	
---------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;
use work.all; 

entity SB_PLL40_2F_PAD_DS  is 
	
	generic ( 
		----------------------------------------------------------------------------------
                --VITAL PARAMETER
                ---------------------------------------------------------------------------------
                TimingChecksOn  	: boolean := true;
                Xon   			: boolean := true;
	        MsgOn 			: boolean := false;
                --- VITAL input port delay 
                tipd_PACKAGEPIN  	: VitalDelayType01 := (0 ns, 0 ns);
                tipd_PACKAGEPINB        : VitalDelayType01 := (0 ns, 0 ns);
            	tipd_EXTFEEDBACK        : VitalDelayType01 := (0 ns, 0 ns);
            	tipd_DYNAMICDELAY       : VitalDelayArrayType01(7 downto 0)  := (others => (0 ns, 0 ns));
            	tipd_BYPASS             : VitalDelayType01 := (0 ns, 0 ns);
            	tipd_RESETB             : VitalDelayType01 := (0 ns, 0 ns);
                tipd_SDI        	: VitalDelayType01 := (0 ns, 0 ns);
            	tipd_SCLK           	: VitalDelayType01 := (0 ns, 0 ns);
            	tipd_LATCHINPUTVALUE   	: VitalDelayType01 := (0 ns, 0 ns);
		-- VITAL Path Delay 	
            	tpd_PACKAGEPIN_PLLOUTCOREA           	: VitalDelayType01 := (0 ns, 0 ns);
            	tpd_PACKAGEPIN_PLLOUTGLOBALA          	: VitalDelayType01 := (0 ns, 0 ns);

            	tpd_PACKAGEPIN_PLLOUTCOREB           	: VitalDelayType01 := (0 ns, 0 ns);
            	tpd_PACKAGEPIN_PLLOUTGLOBALB          	: VitalDelayType01 := (0 ns, 0 ns);
	         -- Entity Parameters 	
		 FEEDBACK_PATH 			: string 		 :="SIMPLE";   -- SIMPLE/DELAY/PHASE_AND_DELAY/EXTERNAL 
		 DELAY_ADJUSTMENT_MODE_FEEDBACK	: string 		 :="FIXED";    -- FIXED/DYNAMIC  
		 DELAY_ADJUSTMENT_MODE_RELATIVE : string 		 :="FIXED";    -- FIXED/DYNAMIC 
		 SHIFTREG_DIV_MODE		: bit_vector(1 downto 0) := "00";      -- 00 (div by 4)/ 01 (div by 7)/11 (div by 5)   	 
		 FDA_FEEDBACK			: bit_vector(3 downto 0) :="0000";
		 FDA_RELATIVE			: bit_vector(3 downto 0) := "0000";
		 PLLOUT_SELECT_PORTA		: string 		 :="GENCLK"; 
		 PLLOUT_SELECT_PORTB		: string 		 :="GENCLK"; 

		 DIVR				: bit_vector(3 downto 0) := "0000";
		 DIVF  				: bit_vector(6 downto 0) := "0000000";
		 DIVQ	   			: bit_vector(2 downto 0) := "000";  
		 FILTER_RANGE 			: bit_vector(2 downto 0) := "000";
		 		
 		 ENABLE_ICEGATE_PORTA	        : bit 			 :='0';
 		 ENABLE_ICEGATE_PORTB	        : bit 			 :='0';
		 TEST_MODE			: bit 			 :='0';  
		 EXTERNAL_DIVIDE_FACTOR         : integer 		 := 1      -- Required for PLL Config Wizard.  
	);
	port (
                PACKAGEPIN		: in std_logic;           -- PLL ref clock(+), driven by PAD.  
                PACKAGEPINB		: in std_logic;           -- PLL ref clock(-), driven by PAD.  
                PLLOUTCOREA	     	: out std_logic;          -- PLLA output to core logic through local routings. 
                PLLOUTGLOBALA           : out std_logic;   	  -- PLLA output to dedicated global clock network
                PLLOUTCOREB	     	: out std_logic;          -- PLLB output to core logic through local routings. 
                PLLOUTGLOBALB           : out std_logic;   	  -- PLLB output to dedicated global clock network
                EXTFEEDBACK             : in std_logic;  	  -- FB driven by core logic
                DYNAMICDELAY            : in std_logic_vector(7 downto 0);  -- driven by core logic
                LOCK                    : out std_logic;	  -- PLL Lock signal output  
                BYPASS                  : in std_logic; 	  -- REFCLK passed to PLLOUT when bypass is '1'.Driven by core logic
                RESETB                  : in std_logic; 	  -- Active low reset,Driven by core logic
                SDI                     : in std_logic;		  -- Test Input. Driven by core logic. 
                SDO                     : out std_logic; 	  -- Test output to RB Logic Tile.
                SCLK                    : in std_logic;	          -- Test Clk input.Driven by core logic. 
                LATCHINPUTVALUE         : in std_logic 		  -- iCEGate signal
	);

       attribute VITAL_LEVEL0 of SB_PLL40_2F_PAD_DS : entity is true;

end SB_PLL40_2F_PAD_DS; 

architecture SB_PLL40_2F_PAD_DS_V of SB_PLL40_2F_PAD_DS is 

	attribute VITAL_LEVEL0 of SB_PLL40_2F_PAD_DS_V  : architecture is true;


 component SbtSPLL40  is
 
	generic ( 
		 FEEDBACK_PATH 			: string 	:="SIMPLE"; 
		 DELAY_ADJUSTMENT_MODE_FEEDBACK	: string 	:="FIXED"; 
		 DELAY_ADJUSTMENT_MODE_RELATIVE : string 	:="FIXED";
		 SHIFTREG_DIV_MODE		: bit_vector(1 downto 0) := "00";	
		 FDA_FEEDBACK			: bit_vector(3 downto 0) :="0000";
		 FDA_RELATIVE			: bit_vector(3 downto 0) := "0000";
		 PLLOUT_SELECT_PORTA		: string 	:="GENCLK"; 
		 PLLOUT_SELECT_PORTB            : string        :="GENCLK"; 

		 DIVR				: bit_vector(3 downto 0) := "0000";
		 DIVF  				: bit_vector(6 downto 0) := "0000000";
		 DIVQ	   			:bit_vector(2 downto 0)  := "000";  
		 FILTER_RANGE 			:bit_vector(2 downto 0)  := "000";
		 		
 		ENABLE_ICEGATE_PORTA             :bit 			:='0';
		ENABLE_ICEGATE_PORTB            :bit 			:='0' 
	);
	port	(
		REFERENCECLK	: in    std_logic;
		EXTFEEDBACK 	: in    std_logic;
		DYNAMICDELAY	: in    std_logic_vector(7 downto 0); 
		BYPASS 		: in	std_logic;
		RESETB	 	: in 	std_logic;
		PLLOUT1 	: out  	std_logic;
		PLLOUT2		: out 	std_logic ; 
		LOCK		: out 	std_logic  
	); 
end component;

  -- Vital Wire Delay Signals   	
  signal PACKAGEPIN_ipd 	: std_ulogic := 'X';
  signal PACKAGEPINB_ipd 	: std_ulogic := 'X';
  signal EXTFEEDBACK_ipd  	: std_ulogic := 'X';
  signal DYNAMICDELAY_ipd  	: std_logic_vector(7 downto 0) := (others =>'X');
  signal BYPASS_ipd   		: std_ulogic := 'X';
  signal RESETB_ipd 		: std_ulogic := 'X';
  signal SDI_ipd  		: std_ulogic := 'X';
  signal SCLK_ipd  		: std_ulogic := 'X';
  signal LATCHINPUTVALUE_ipd  	: std_ulogic := 'X';

 -- Vital output logic signals
 signal PLLOUTCOREA_zd : std_ulogic;
 signal PLLOUTGLOBALA_zd : std_ulogic;
 signal PLLOUTCOREB_zd : std_ulogic;
 signal PLLOUTGLOBALB_zd : std_ulogic;
 signal LOCK_zd : std_ulogic;
 signal SDO_zd : std_ulogic;
 signal Violation : std_ulogic;

 -- Functional signals 
 signal not_resetb  		 : std_logic; 
 signal SPLLOUT1net, SPLLOUT2net : std_logic; 
 signal PLLOUTCOREA_temp 	 : std_logic; 
 signal PLLOUTGLOBALA_temp 	 : std_logic; 
 signal PLLOUTCOREB_temp 	 : std_logic; 
 signal PLLOUTGLOBALB_temp 	 : std_logic; 


begin 

 WireDelay   : block
 begin
          VitalWireDelay (PACKAGEPIN_ipd, PACKAGEPIN, tipd_PACKAGEPIN);
          VitalWireDelay (PACKAGEPINB_ipd, PACKAGEPINB, tipd_PACKAGEPINB);
          VitalWireDelay (EXTFEEDBACK_ipd,  EXTFEEDBACK, tipd_EXTFEEDBACK);
	  DYNAMIC_DELAY : for i in 7 downto 0 generate 
	          VitalWireDelay (DYNAMICDELAY_ipd(i),DYNAMICDELAY(i),tipd_DYNAMICDELAY(i));
	  end generate DYNAMIC_DELAY; 
          VitalWireDelay (BYPASS_ipd,BYPASS, tipd_BYPASS);
          VitalWireDelay (RESETB_ipd,RESETB, tipd_RESETB);
          VitalWireDelay (SDI_ipd, SDI, tipd_SDI);
          VitalWireDelay (SCLK_ipd, SCLK, tipd_SCLK);
          VitalWireDelay (LATCHINPUTVALUE_ipd, LATCHINPUTVALUE, tipd_LATCHINPUTVALUE);
 end block;

 ------ Behavioral Section   
 not_resetb <= not(RESETB_ipd);  

 instSbtSPLL : SbtSPLL40 
 generic map 	( 
		FEEDBACK_PATH 			=> FEEDBACK_PATH,
		DELAY_ADJUSTMENT_MODE_RELATIVE 	=> DELAY_ADJUSTMENT_MODE_RELATIVE,
		DELAY_ADJUSTMENT_MODE_FEEDBACK 	=> DELAY_ADJUSTMENT_MODE_FEEDBACK,
		SHIFTREG_DIV_MODE 		=> SHIFTREG_DIV_MODE,
		FDA_RELATIVE 			=> FDA_RELATIVE,
		FDA_FEEDBACK 			=> FDA_FEEDBACK,
		PLLOUT_SELECT_PORTA 		=> PLLOUT_SELECT_PORTA,
		PLLOUT_SELECT_PORTB 		=> PLLOUT_SELECT_PORTB, 
		DIVR 				=> DIVR,
		DIVF 				=> DIVF,
		DIVQ 				=> DIVQ,
		FILTER_RANGE 			=> FILTER_RANGE,
 		ENABLE_ICEGATE_PORTA             =>'0',
		ENABLE_ICEGATE_PORTB            =>'0' 
	     	)
 port map    	(
                REFERENCECLK 			=> PACKAGEPIN_ipd,
                EXTFEEDBACK 			=> EXTFEEDBACK_ipd,
                DYNAMICDELAY 			=> DYNAMICDELAY_ipd,
                BYPASS 				=> BYPASS_ipd,
                RESETB 				=> not_resetb ,
                PLLOUT1 			=> SPLLOUT1net,
                PLLOUT2 			=> SPLLOUT2net,
                LOCK 				=> LOCK
		);


  -- PLLA
 process(PLLOUTCOREA_temp, SPLLOUT1net)  
 begin 
	if(ENABLE_ICEGATE_PORTA = '1' and LATCHINPUTVALUE_ipd ='1') then 
		PLLOUTCOREA_temp <= PLLOUTCOREA_temp ; 
	else 
		PLLOUTCOREA_temp <= SPLLOUT1net; 
	end if;
 end process; 


 process(PLLOUTGLOBALA_temp, SPLLOUT1net)  
 begin 
	if(ENABLE_ICEGATE_PORTA = '1' and LATCHINPUTVALUE_ipd ='1') then 
		PLLOUTGLOBALA_temp <= PLLOUTGLOBALA_temp ; 
	else 
		PLLOUTGLOBALA_temp <= SPLLOUT1net; 
	end if; 
 end process; 

 PLLOUTCOREA_zd 	<= PLLOUTCOREA_temp; 
 PLLOUTGLOBALA_zd 	<= PLLOUTGLOBALA_temp;  

 --PLLB

 process(PLLOUTCOREB_temp, SPLLOUT2net)  
 begin 
	if(ENABLE_ICEGATE_PORTB = '1' and LATCHINPUTVALUE_ipd ='1') then 
		PLLOUTCOREB_temp <= PLLOUTCOREB_temp ; 
	else 
		PLLOUTCOREB_temp <= SPLLOUT2net; 
	end if;
 end process; 


 process(PLLOUTGLOBALB_temp, SPLLOUT2net)  
 begin 
	if(ENABLE_ICEGATE_PORTB = '1' and LATCHINPUTVALUE_ipd ='1') then 
		PLLOUTGLOBALB_temp <= PLLOUTGLOBALB_temp ; 
	else 
		PLLOUTGLOBALB_temp <= SPLLOUT2net; 
	end if; 
 end process; 

 PLLOUTCOREB_zd 	<= PLLOUTCOREB_temp; 
 PLLOUTGLOBALB_zd 	<= PLLOUTGLOBALB_temp;  
 
 ---------------------------- 
 -- Vital Path delay  
 ---------------------------
  VITALPathDelay          : process (PLLOUTCOREA_zd, PLLOUTGLOBALA_zd,PLLOUTCOREB_zd, PLLOUTGLOBALB_zd,PACKAGEPIN_ipd )
  	variable PLLOUTCOREA_GlitchData 	: VitalGlitchDataType;
	variable PLLOUTGLOBALA_GlitchData 	: VitalGlitchDataType;
  	variable PLLOUTCOREB_GlitchData 	: VitalGlitchDataType;
	variable PLLOUTGLOBALB_GlitchData 	: VitalGlitchDataType;
	variable LOCK_zd		 	: VitalGlitchDataType;

  begin 		
  VitalPathDelay01 (
      OutSignal                 => PLLOUTCOREA,
      GlitchData                => PLLOUTCOREA_GlitchData,
      OutSignalName             => "PLLOUTCOREA",
      OutTemp                   => PLLOUTCOREA_zd,
      Paths                     => (0 => (PACKAGEPIN_ipd'last_event, tpd_PACKAGEPIN_PLLOUTCOREA,true)
							),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
	  
  VitalPathDelay01 (
      OutSignal                 => PLLOUTGLOBALA,
      GlitchData                => PLLOUTGLOBALA_GlitchData,
      OutSignalName             => "PLLOUTGLOBALA",
      OutTemp                   => PLLOUTGLOBALA_zd,
      Paths                     => (0 => (PACKAGEPIN_ipd'last_event, tpd_PACKAGEPIN_PLLOUTGLOBALA, true)
									),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

  VitalPathDelay01 (
      OutSignal                 => PLLOUTCOREB,
      GlitchData                => PLLOUTCOREB_GlitchData,
      OutSignalName             => "PLLOUTCOREB",
      OutTemp                   => PLLOUTCOREB_zd,
      Paths                     => (0 => (PACKAGEPIN_ipd'last_event, tpd_PACKAGEPIN_PLLOUTCOREB,true)
							),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
	  
  VitalPathDelay01 (
      OutSignal                 => PLLOUTGLOBALB,
      GlitchData                => PLLOUTGLOBALB_GlitchData,
      OutSignalName             => "PLLOUTGLOBALB",
      OutTemp                   => PLLOUTGLOBALB_zd,
      Paths                     => (0 => (PACKAGEPIN_ipd'last_event, tpd_PACKAGEPIN_PLLOUTGLOBALB, true)
									),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
 end process VITALPathDelay;	

end SB_PLL40_2F_PAD_DS_V; 


---------------------------------------------------------------------------
----		 	SB_TMDS_deserilizer(HDMI)			---	
---------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;

entity SB_TMDS_deserializer is 
	generic 	(
	----------------------------------------------------------------------------------
        --VITAL PARAMETER
	---------------------------------------------------------------------------------
	TimingChecksOn  	: boolean := true;
	Xon   			: boolean := true;
	MsgOn 			: boolean := true;
	--- VITAL input port delay 
	tipd_TMDSch0p	  			: VitalDelayType01 := (0 ns, 0 ns);
	tipd_TMDSch0n  				: VitalDelayType01 := (0 ns, 0 ns);
	tipd_TMDSch1p 	       			: VitalDelayType01 := (0 ns, 0 ns);
	tipd_TMDSch1n 	       			: VitalDelayType01 := (0 ns, 0 ns);
	tipd_TMDSch2p 	       			: VitalDelayType01 := (0 ns, 0 ns);
	tipd_TMDSch2n 	       			: VitalDelayType01 := (0 ns, 0 ns);
	tipd_TMDSclkp 	       			: VitalDelayType01 := (0 ns, 0 ns);
	tipd_TMDSclkn 	       			: VitalDelayType01 := (0 ns, 0 ns);
	tipd_RSTNdeser 	       			: VitalDelayType01 := (0 ns, 0 ns);
	tipd_RSTNpll	       			: VitalDelayType01 := (0 ns, 0 ns);
	tipd_EN	       				: VitalDelayType01 := (0 ns, 0 ns);
	tipd_PHASELch0 	       			: VitalDelayArrayType01( 3 downto 0 )  :=(others => (0 ns, 0 ns));
	tipd_PHASELch1 	       			: VitalDelayArrayType01( 3 downto 0 )  :=(others => (0 ns, 0 ns)); 
	tipd_PHASELch2 	       			: VitalDelayArrayType01( 3 downto 0 )  :=(others => (0 ns, 0 ns)); 
	tipd_EXTFEEDBACK       			: VitalDelayType01 := (0 ns, 0 ns);
	tipd_DYNAMICDELAY       		: VitalDelayArrayType01( 7 downto 0 )  :=(others => (0 ns, 0 ns));
	tipd_BYPASS 	       			: VitalDelayType01 := (0 ns, 0 ns);
	tipd_LATCHINPUTVALUE 	       		: VitalDelayType01 := (0 ns, 0 ns);
	tipd_SDI       				: VitalDelayType01 := (0 ns, 0 ns);
	tipd_SCLK	       			: VitalDelayType01 := (0 ns, 0 ns);
	-- VITAL Path Delay 	
	tpd_TMDSclkp_PLLOUTGLOBALclkx1         	: VitalDelayType01 := (0 ns, 0 ns);
	tpd_TMDSclkp_PLLOUTCOREclkx1 	     	: VitalDelayType01 := (0 ns, 0 ns);
	tpd_TMDSclkp_PLLOUTGLOBALclkx5         	: VitalDelayType01 := (0 ns, 0 ns);
	tpd_TMDSclkp_PLLOUTCOREclkx5           	: VitalDelayType01 := (0 ns, 0 ns);
	-- VITAL clk-to-output path delay
        tpd_TMDSclkp_RAWDATAch0_posedge 	: VitalDelayArrayType01( 9 downto 0) := (others => (0 ns, 0 ns));
        tpd_TMDSclkp_RAWDATAch1_posedge 	: VitalDelayArrayType01( 9 downto 0) := (others => (0 ns, 0 ns));
        tpd_TMDSclkp_RAWDATAch2_posedge 	: VitalDelayArrayType01( 9 downto 0) := (others => (0 ns, 0 ns));
	-- VITAL Setup delays 
        tsetup_TMDSch0p_TMDSclkp_posedge_posedge 		: VitalDelayType                   := 0 ns; 
   	tsetup_TMDSch0p_TMDSclkp_negedge_posedge	 	: VitalDelayType                   := 0 ns; 
        tsetup_TMDSch0p_TMDSclkp_posedge_negedge 		: VitalDelayType                   := 0 ns; 
   	tsetup_TMDSch0p_TMDSclkp_negedge_negedge	 	: VitalDelayType                   := 0 ns; 
        tsetup_TMDSch0n_TMDSclkp_posedge_posedge 		: VitalDelayType                   := 0 ns; 
   	tsetup_TMDSch0n_TMDSclkp_negedge_posedge	 	: VitalDelayType                   := 0 ns; 
        tsetup_TMDSch0n_TMDSclkp_posedge_negedge 		: VitalDelayType                   := 0 ns; 
   	tsetup_TMDSch0n_TMDSclkp_negedge_negedge	 	: VitalDelayType                   := 0 ns; 

        tsetup_TMDSch1p_TMDSclkp_posedge_posedge 		: VitalDelayType                   := 0 ns; 
   	tsetup_TMDSch1p_TMDSclkp_negedge_posedge	 	: VitalDelayType                   := 0 ns; 
        tsetup_TMDSch1p_TMDSclkp_posedge_negedge 		: VitalDelayType                   := 0 ns; 
   	tsetup_TMDSch1p_TMDSclkp_negedge_negedge	 	: VitalDelayType                   := 0 ns; 
        tsetup_TMDSch1n_TMDSclkp_posedge_posedge 		: VitalDelayType                   := 0 ns; 
   	tsetup_TMDSch1n_TMDSclkp_negedge_posedge	 	: VitalDelayType                   := 0 ns; 
        tsetup_TMDSch1n_TMDSclkp_posedge_negedge 		: VitalDelayType                   := 0 ns; 
   	tsetup_TMDSch1n_TMDSclkp_negedge_negedge	 	: VitalDelayType                   := 0 ns; 

        tsetup_TMDSch2p_TMDSclkp_posedge_posedge 		: VitalDelayType                   := 0 ns; 
   	tsetup_TMDSch2p_TMDSclkp_negedge_posedge	 	: VitalDelayType                   := 0 ns; 
        tsetup_TMDSch2p_TMDSclkp_posedge_negedge 		: VitalDelayType                   := 0 ns; 
   	tsetup_TMDSch2p_TMDSclkp_negedge_negedge	 	: VitalDelayType                   := 0 ns; 
        tsetup_TMDSch2n_TMDSclkp_posedge_posedge 		: VitalDelayType                   := 0 ns; 
   	tsetup_TMDSch2n_TMDSclkp_negedge_posedge	 	: VitalDelayType                   := 0 ns; 
        tsetup_TMDSch2n_TMDSclkp_posedge_negedge 		: VitalDelayType                   := 0 ns; 
   	tsetup_TMDSch2n_TMDSclkp_negedge_negedge	 	: VitalDelayType                   := 0 ns; 

	-- VITAL Hold delays 
        thold_TMDSch0p_TMDSclkp_posedge_posedge 		: VitalDelayType                   := 0 ns; 
   	thold_TMDSch0p_TMDSclkp_negedge_posedge	 		: VitalDelayType                   := 0 ns; 
        thold_TMDSch0p_TMDSclkp_posedge_negedge 		: VitalDelayType                   := 0 ns; 
        thold_TMDSch0p_TMDSclkp_negedge_negedge 		: VitalDelayType                   := 0 ns; 
        thold_TMDSch0n_TMDSclkp_posedge_posedge 		: VitalDelayType                   := 0 ns; 
   	thold_TMDSch0n_TMDSclkp_negedge_posedge	 		: VitalDelayType                   := 0 ns; 
        thold_TMDSch0n_TMDSclkp_posedge_negedge 		: VitalDelayType                   := 0 ns; 
        thold_TMDSch0n_TMDSclkp_negedge_negedge 		: VitalDelayType                   := 0 ns; 

        thold_TMDSch1p_TMDSclkp_posedge_posedge 		: VitalDelayType                   := 0 ns; 
   	thold_TMDSch1p_TMDSclkp_negedge_posedge	 		: VitalDelayType                   := 0 ns; 
        thold_TMDSch1p_TMDSclkp_posedge_negedge 		: VitalDelayType                   := 0 ns; 
        thold_TMDSch1p_TMDSclkp_negedge_negedge 		: VitalDelayType                   := 0 ns; 
        thold_TMDSch1n_TMDSclkp_posedge_posedge 		: VitalDelayType                   := 0 ns; 
   	thold_TMDSch1n_TMDSclkp_negedge_posedge	 		: VitalDelayType                   := 0 ns; 
        thold_TMDSch1n_TMDSclkp_posedge_negedge 		: VitalDelayType                   := 0 ns; 
        thold_TMDSch1n_TMDSclkp_negedge_negedge 		: VitalDelayType                   := 0 ns; 

        thold_TMDSch2p_TMDSclkp_posedge_posedge 		: VitalDelayType                   := 0 ns; 
   	thold_TMDSch2p_TMDSclkp_negedge_posedge	 		: VitalDelayType                   := 0 ns; 
        thold_TMDSch2p_TMDSclkp_posedge_negedge 		: VitalDelayType                   := 0 ns; 
        thold_TMDSch2p_TMDSclkp_negedge_negedge 		: VitalDelayType                   := 0 ns; 
        thold_TMDSch2n_TMDSclkp_posedge_posedge 		: VitalDelayType                   := 0 ns; 
   	thold_TMDSch2n_TMDSclkp_negedge_posedge	 		: VitalDelayType                   := 0 ns; 
        thold_TMDSch2n_TMDSclkp_posedge_negedge 		: VitalDelayType                   := 0 ns; 
        thold_TMDSch2n_TMDSclkp_negedge_negedge 		: VitalDelayType                   := 0 ns; 
	--- DVI generic params 
	 FEEDBACK_PATH 			: string 		:= "PHASE_AND_DELAY" ;	   
	 DELAY_ADJUSTMENT_MODE_FEEDBACK : string 		:= "FIXED"; 
	 DELAY_ADJUSTMENT_MODE_RELATIVE : string		:= "FIXED"; 
	 SHIFTREG_DIV_MODE		: bit_vector(1 downto 0):= "11"; 		--Set to div by 5 mode 
	 FDA_FEEDBACK			: bit_vector(3 downto 0):="0000"; 		
	 FDA_RELATIVE 			: bit_vector(3 downto 0):= "0000";  
	 PLLOUT_SELECT_PORTA 		: string 		:= "GENCLK";    	-- Clkx5
	 PLLOUT_SELECT_PORTB 		: string 		:= "SHIFTREG_0deg"; 	-- Clkx1
	-- Frequency Parameters: Current defaults are for TMDS Clk = 30-40MHz 
	 DIVR 				: bit_vector(3 downto 0) := "0000"; 	
	 DIVF 				: bit_vector(6 downto 0) := "0000000"; 
	 DIVQ 				: bit_vector(2 downto 0) := "010"; 	
	 FILTER_RANGE 			: bit_vector(2 downto 0) := "011"; 	
	 ENABLE_ICEGATE_PORTA 		: bit			 := '0';
	 ENABLE_ICEGATE_PORTB 		: bit 			 := '0';
	-- Test Mode parameter
	 TEST_MODE 			: bit 			 := '0';
	 EXTERNAL_DIVIDE_FACTOR 	: integer		  := 1 		-- Required for  PLL Config Wizard.
	); 
	port	( 
        -- TMDS input interface
  	TMDSch0p		: in 	std_logic ;             		-- TMDS ch 0 differential input pos
	TMDSch0n		: in	std_logic ;             		-- TMDS ch 0 differential input neg
	TMDSch1p		: in	std_logic ; 	          		-- TMDS ch 1 differential input pos
	TMDSch1n		: in	std_logic ;   	        		-- TMDS ch 1 differential input neg
   	TMDSch2p		: in	std_logic ; 	        		-- TMDS ch 2 differential input pos
   	TMDSch2n		: in 	std_logic ;             		-- TMDS ch 2 differential input neg
   	TMDSclkp		: in	std_logic ;             		-- TMDS clock differential input pos
   	TMDSclkn		: in	std_logic ;             		-- TMDS clock differential input neg                                
        -- Receiver controller interface
  	RSTNdeser		: in 	std_logic ;             		-- Reset deserailzier logics- active low
	RSTNpll			: in	std_logic ;             		-- Reset deserializer PLL- active low
   	EN			: in	std_logic ;             		-- Enable deserializer- active high
    	PHASELch0		: in	std_logic_vector( 3 downto 0) ; 	--  Clock phase delay compensation select for ch 0
   	PHASELch1		: in	std_logic_vector( 3 downto 0) ; 	--  Clock phase delay compensation select for ch 1
   	PHASELch2		: in	std_logic_vector( 3 downto 0) ; 	--  Clock phase delay compensation select for ch 2
   	PLLlock			: out 	std_logic ;              	 	--  PLL lock signal- active high
   	PLLOUTGLOBALclkx1 	: out 	std_logic ;     			--  PLL output on global n/w 
   	PLLOUTCOREclkx1 	: out 	std_logic ;      			--  PLL output on global n/w 
   	PLLOUTGLOBALclkx5 	: out 	std_logic ; 	 			--  PLL output on global n/w 
   	PLLOUTCOREclkx5 	: out 	std_logic ;      			--  PLL output on global n/w
   	RAWDATAch0 		: out 	std_logic_vector( 9 downto 0) ;     	--  Recovered ch 0 10-bit data 
   	RAWDATAch1 		: out	std_logic_vector( 9 downto 0) ;     	--  Recovered ch 1 10-bit data
   	RAWDATAch2 		: out 	std_logic_vector( 9 downto 0) ;     	--  Recovered ch 2 10-bit data
  	EXTFEEDBACK	  	: in 	std_logic ;   			    	--  Driven by core logic. Not required HDMI mode.
  	DYNAMICDELAY 		: in 	std_logic_vector ( 7 downto 0 ) ;   	--  Driven by core logic. Not required for HDMI mode.
  	BYPASS			: in 	std_logic ; 		    		--  Driven by core logic. Not required for HDMI mode.
  	LATCHINPUTVALUE 	: in 	std_logic ;  		    		--  iCEGate signal. Not required for HDMI mode
	-- Test Pins
  	SDO 			: out 	std_logic ; 		    		--  Output of PLL
  	SDI			: in 	std_logic ; 		    		--  Driven by core logic
  	SCLK			: in    std_logic 		    		--  Driven by core logic
  	);


	attribute VITAL_LEVEL0 of SB_TMDS_deserializer : entity is true;

end  SB_TMDS_deserializer;  

architecture SB_TMDS_deserializer_V  of SB_TMDS_deserializer is 

  attribute VITAL_LEVEL0 of SB_TMDS_deserializer_V : architecture is true;

  component dvi_deserializer is
  	port ( 
		en  	: in 	std_logic ; 							
		rstn  	: in 	std_logic ; 
		din		: in	std_logic ; 
		clkx5in	: in	std_logic ; 	
		clkx1in	: in 	std_logic ; 
		rawdata : out  	std_logic_vector(9 downto 0)	
	      ); 	
  end component ; 
  
  component clkdelay16 is 
	generic (
		BUF_DELAY : time  		:= 100 ps  
		); 		
	port    ( 
		dlyin    : in 	 	std_logic;  
		dlyout	 : out 		std_logic ;  
		dly_sel	 : in 		std_logic_vector( 3 downto 0)
		); 															  	
  end component;
  
  component  SB_PLL40_2F_PAD_DS  is 	
	generic ( 
	----------------------------------------------------------------------------------
        --VITAL PARAMETER
        ---------------------------------------------------------------------------------
        TimingChecksOn  	: boolean := true;
        Xon   			: boolean := true;
    	MsgOn 			: boolean := false;
        --- VITAL input port delay 
        tipd_PACKAGEPIN  	: VitalDelayType01 := (0 ns, 0 ns);
        tipd_PACKAGEPINB        : VitalDelayType01 := (0 ns, 0 ns);
        tipd_EXTFEEDBACK        : VitalDelayType01 := (0 ns, 0 ns);
        tipd_DYNAMICDELAY       : VitalDelayArrayType01(7 downto 0)  := (others => (0 ns, 0 ns));
        tipd_BYPASS             : VitalDelayType01 := (0 ns, 0 ns);
        tipd_RESETB             : VitalDelayType01 := (0 ns, 0 ns);
        tipd_SDI        	: VitalDelayType01 := (0 ns, 0 ns);
        tipd_SCLK           	: VitalDelayType01 := (0 ns, 0 ns);
        tipd_LATCHINPUTVALUE   	: VitalDelayType01 := (0 ns, 0 ns);
		-- VITAL Path Delay 	
        tpd_PACKAGEPIN_PLLOUTCOREA           	: VitalDelayType01 := (0 ns, 0 ns);
        tpd_PACKAGEPIN_PLLOUTGLOBALA          	: VitalDelayType01 := (0 ns, 0 ns);

        tpd_PACKAGEPIN_PLLOUTCOREB           	: VitalDelayType01 := (0 ns, 0 ns);
        tpd_PACKAGEPIN_PLLOUTGLOBALB          	: VitalDelayType01 := (0 ns, 0 ns);
	     -- Entity Parameters 	
	FEEDBACK_PATH 				: string 		 :="SIMPLE";   -- SIMPLE/DELAY/PHASE_AND_DELAY/EXTERNAL 
	DELAY_ADJUSTMENT_MODE_FEEDBACK		: string 		 :="FIXED";    -- FIXED/DYNAMIC  
	DELAY_ADJUSTMENT_MODE_RELATIVE 		: string 		 :="FIXED";    -- FIXED/DYNAMIC 
	SHIFTREG_DIV_MODE			: bit_vector(1 downto 0) := "11";      -- 00 (div by 4)/ 01 (div by 7)/11 (div by 5)   	 
	FDA_FEEDBACK				: bit_vector(3 downto 0) :="0000";
	FDA_RELATIVE				: bit_vector(3 downto 0) := "0000";
	PLLOUT_SELECT_PORTA			: string 		 :="GENCLK"; 
	PLLOUT_SELECT_PORTB			: string 		 :="GENCLK"; 

	DIVR					: bit_vector(3 downto 0) := "0000";
	DIVF  					: bit_vector(6 downto 0) := "0000000";
	DIVQ	   				: bit_vector(2 downto 0) := "000";  
	FILTER_RANGE 				: bit_vector(2 downto 0) := "000";
	 		
 	ENABLE_ICEGATE_PORTA			: bit 			 :='0';
 	ENABLE_ICEGATE_PORTB			: bit 			 :='0';
	TEST_MODE				: bit 			 :='0';  
	EXTERNAL_DIVIDE_FACTOR         		: integer 		 := 1      -- Required for PLL Config Wizard.  
	);
	port (
        PACKAGEPIN				: in std_logic;           -- PLL ref clock(+), driven by PAD.  
        PACKAGEPINB				: in std_logic;           -- PLL ref clock(-), driven by PAD.  
        PLLOUTCOREA	     			: out std_logic;          -- PLLA output to core logic through local routings. 
        PLLOUTGLOBALA           		: out std_logic;   	  	  -- PLLA output to dedicated global clock network
        PLLOUTCOREB	     			: out std_logic;          -- PLLB output to core logic through local routings. 
        PLLOUTGLOBALB           		: out std_logic;   	  -- PLLB output to dedicated global clock network
        EXTFEEDBACK             		: in std_logic;  	  -- FB driven by core logic
        DYNAMICDELAY            		: in std_logic_vector(7 downto 0);  -- driven by core logic
        LOCK                    		: out std_logic;	  -- PLL Lock signal output  
        BYPASS                  		: in std_logic; 	  -- REFCLK passed to PLLOUT when bypass is '1'.Driven by core logic
        RESETB                  		: in std_logic; 	  -- Active low reset,Driven by core logic
        SDI                     		: in std_logic;		  -- Test Input. Driven by core logic. 
        SDO                     		: out std_logic; 	  -- Test output to RB Logic Tile.
        SCLK                    		: in std_logic;	          -- Test Clk input.Driven by core logic. 
        LATCHINPUTVALUE         		: in std_logic 		  -- iCEGate signal
	);	
end component;

	signal clk1xout_global, clk5xout_global 	: std_logic ;  
    	signal clk1xout_core, clk5xout_core		: std_logic ; 
  
  	signal ch0_clk5xin	: std_logic ; 
  	signal ch1_clk5xin	: std_logic ; 
  	signal ch2_clk5xin	: std_logic ; 	
        --- Vital Signals 
	signal  TMDSch0p_ipd	      : std_ulogic := 'X';
        signal  TMDSch0n_ipd	      : std_ulogic := 'X';
        signal  TMDSch1p_ipd          : std_ulogic := 'X';
        signal  TMDSch1n_ipd          : std_ulogic := 'X';
        signal  TMDSch2p_ipd          : std_ulogic := 'X';
        signal  TMDSch2n_ipd          : std_ulogic := 'X';
        signal  TMDSclkp_ipd          : std_ulogic := 'X';
        signal  TMDSclkn_ipd          : std_ulogic := 'X';
        signal  RSTNdeser_ipd         : std_ulogic := 'X';
        signal  RSTNpll_ipd           : std_ulogic := 'X';
        signal  EN_ipd      	      : std_ulogic := 'X';
        signal  PHASELch0_ipd         : std_logic_vector( 3 downto 0) := (others => 'X');
        signal  PHASELch1_ipd         : std_logic_vector( 3 downto 0) := (others => 'X');
        signal  PHASELch2_ipd         : std_logic_vector( 3 downto 0) := (others => 'X');
        signal  EXTFEEDBACK_ipd       : std_ulogic := 'X';
        signal  DYNAMICDELAY_ipd      : std_logic_vector(7 downto 0) := (others => 'X');
        signal  BYPASS_ipd            : std_ulogic := 'X'; 
        signal  LATCHINPUTVALUE_ipd   : std_ulogic := 'X'; 
        signal  SDI_ipd               : std_ulogic := 'X'; 
        signal  SCLK_ipd              : std_ulogic := 'X'; 

	signal  RAWDATAch0_zd 	      : std_logic_vector( 9 downto 0); 
	signal  RAWDATAch1_zd 	      : std_logic_vector( 9 downto 0); 
	signal  RAWDATAch2_zd 	      : std_logic_vector( 9 downto 0); 
	signal	PLLOUTGLOBALclkx1_zd  : std_ulogic ; 
	signal	PLLOUTCOREclkx1_zd    : std_ulogic ; 
	signal 	PLLOUTGLOBALclkx5_zd  : std_ulogic ;
	signal  PLLOUTCOREclkx5_zd    : std_ulogic ; 
	signal  PLLlock_zd	      : std_ulogic ;
	signal	SDO_zd	     	      : std_ulogic ;
     				
begin 

 WireDelay   : block
 begin
          VitalWireDelay (TMDSch0p_ipd,TMDSch0p, tipd_TMDSch0p );
          VitalWireDelay (TMDSch0n_ipd,TMDSch0n, tipd_TMDSch0n );
          VitalWireDelay (TMDSch1p_ipd,TMDSch1p, tipd_TMDSch1p );
          VitalWireDelay (TMDSch1n_ipd,TMDSch1n, tipd_TMDSch1n );
          VitalWireDelay (TMDSch2p_ipd,TMDSch2p, tipd_TMDSch2p );
          VitalWireDelay (TMDSch2n_ipd,TMDSch2n, tipd_TMDSch2n );
          VitalWireDelay (TMDSclkp_ipd,TMDSclkp, tipd_TMDSclkp );
          VitalWireDelay (TMDSclkn_ipd,TMDSclkn, tipd_TMDSclkn );
          VitalWireDelay (RSTNdeser_ipd , RSTNdeser, tipd_RSTNdeser );
	  VitalWireDelay (RSTNpll_ipd, RSTNpll, tipd_RSTNpll ); 
	  VitalWireDelay (EN_ipd, EN, tipd_EN ); 
	  PHASEADJ_DELAY : for i in 3 downto 0 generate
      	    VitalWireDelay (PHASELch0_ipd(i), PHASELch0(i), tipd_PHASELch0(i));
      	    VitalWireDelay (PHASELch1_ipd(i), PHASELch1(i), tipd_PHASELch1(i));
      	    VitalWireDelay (PHASELch2_ipd(i), PHASELch2(i), tipd_PHASELch2(i));
    	  end generate PHASEADJ_DELAY ;
	  VitalWireDelay (EXTFEEDBACK_ipd, EXTFEEDBACK, tipd_EXTFEEDBACK ); 
	  DYNAMIC_DELAY : for i in 7 downto 0 generate
      	    VitalWireDelay (DYNAMICDELAY_ipd(i), DYNAMICDELAY(i), tipd_DYNAMICDELAY(i));
    	  end generate DYNAMIC_DELAY ;
	  VitalWireDelay (BYPASS_ipd, BYPASS, tipd_BYPASS ); 
	  VitalWireDelay (LATCHINPUTVALUE_ipd , LATCHINPUTVALUE, tipd_LATCHINPUTVALUE ); 
	  VitalWireDelay (SDI_ipd, SDI, tipd_SDI  ); 
	  VitalWireDelay (SCLK_ipd , SCLK, tipd_SCLK  ); 
 end block;

	-- Behavioral  section 
	dviPLL_i : SB_PLL40_2F_PAD_DS  
		generic map (  
		FEEDBACK_PATH				=> "PHASE_AND_DELAY" , 
		DELAY_ADJUSTMENT_MODE_FEEDBACK  	=> "FIXED" ,
		FDA_FEEDBACK 				=> "0000" , 
		DELAY_ADJUSTMENT_MODE_RELATIVE 		=> "FIXED" , 
		FDA_RELATIVE 				=> "0000" , 
		SHIFTREG_DIV_MODE			=> "11" ,
		PLLOUT_SELECT_PORTA			=> "GENCLK" ,
		PLLOUT_SELECT_PORTB			=> "SHIFTREG_0deg" , 
		ENABLE_ICEGATE_PORTA			=> '0' ,
		ENABLE_ICEGATE_PORTB			=> '0' ,
		DIVR					=> "0000" ,   	   	  -- 1  
		DIVF					=> "0000000" ,     	  -- 1
		DIVQ					=> "010" , 		      --Divide VCO out by 2^2 = 4 ; 
		FILTER_RANGE 				=> "011"     
		) 											  	
		port map (	
		PACKAGEPIN 		=> TMDSclkp_ipd ,
            	PACKAGEPINB		=> TMDSclkn_ipd ,
		PLLOUTCOREA 		=> clk5xout_core ,
            	PLLOUTCOREB 		=> clk1xout_core ,
            	PLLOUTGLOBALA 		=> clk5xout_global ,
            	PLLOUTGLOBALB 		=> clk1xout_global ,
            	EXTFEEDBACK	  	=> EXTFEEDBACK_ipd ,
            	DYNAMICDELAY		=> DYNAMICDELAY_ipd ,
            	RESETB			=> RSTNpll_ipd ,
            	BYPASS			=> '0',
            	LATCHINPUTVALUE		=> '0', 
            	LOCK			=> PLLlock,
            	SDI			=> SDI_ipd , 
            	SDO			=> SDO, 
            	SCLK			=> SCLK_ipd
		);
		
	-----------------------------------------------
	PLLOUTGLOBALclkx1_zd <=  clk1xout_global ;  
	PLLOUTCOREclkx1_zd   <=  clk1xout_core; 
	PLLOUTGLOBALclkx5_zd <=  clk5xout_global; 
	PLLOUTCOREclkx5_zd   <=  clk5xout_core; 
	
	 -- channel 0  	
	clkdelay16_ch0_i: clkdelay16
		port map (
			dlyin	=> clk5xout_global, 
			dlyout	=> ch0_clk5xin, 
			dly_sel	=> PHASELch0_ipd 
			);
	
	deserializer_ch0_i : dvi_deserializer 
		port map (
			en	=> EN_ipd,							
			rstn	=> RSTNdeser_ipd, 	 
			din	=> TMDSch0p_ipd	, 
			clkx5in	=> ch0_clk5xin,	
			clkx1in => TMDSclkp_ipd,
			rawdata => RAWDATAch0_zd 
			); 
	-- channel 1 	
	clkdelay16_ch1_i : clkdelay16 
		port map (
			dlyin	=> clk5xout_global, 
			dlyout	=> ch1_clk5xin, 
			dly_sel	=> PHASELch1_ipd 
			);								
	
	deserializer_ch1_i : dvi_deserializer 
		port map (
			en 	=> EN_ipd,							
			rstn	=> RSTNdeser_ipd, 	 
			din	=> TMDSch1p_ipd, 
			clkx5in	=> ch1_clk5xin,	
			clkx1in	=> TMDSclkp_ipd,
			rawdata => RAWDATAch1_zd 
			); 	
	-- Channel 2 
	clkdelay16_ch2_i: clkdelay16 
		port map (
			dlyin 	=> clk5xout_global, 
			dlyout 	=> ch2_clk5xin, 
			dly_sel	=> PHASELch2_ipd 
			);		
	deserializer_ch2_i: dvi_deserializer 
		port map (
			en 	=> EN_ipd,							
			rstn 	=> RSTNdeser_ipd, 	 
			din	=> TMDSch2p_ipd, 
			clkx5in	=> ch2_clk5xin,	
			clkx1in	=> TMDSclkp_ipd,
			rawdata	=> RAWDATAch2_zd 
			); 	

-------------------------------------------------------------------
--VITAL timing check
------------------------------------------------------------------
  VITALTimingCheck : process (TMDSch0p_ipd,TMDSch0n_ipd, TMDSch1p_ipd, TMDSch1n_ipd, TMDSch2p_ipd, TMDSch2n_ipd, TMDSclkp_ipd)
        variable Tviol_TMDSch0p_TMDSclkp_posedge       	: std_ulogic := '0';
        variable Tviol_TMDSch0p_TMDSclkp_negedge 	: std_ulogic := '0';
        variable Tviol_TMDSch0n_TMDSclkp_posedge     	: std_ulogic := '0';
        variable Tviol_TMDSch0n_TMDSclkp_negedge        : std_ulogic := '0';
        variable Tviol_TMDSch1p_TMDSclkp_posedge       	: std_ulogic := '0';
        variable Tviol_TMDSch1p_TMDSclkp_negedge 	: std_ulogic := '0';
        variable Tviol_TMDSch1n_TMDSclkp_posedge     	: std_ulogic := '0';
        variable Tviol_TMDSch1n_TMDSclkp_negedge        : std_ulogic := '0';
        variable Tviol_TMDSch2p_TMDSclkp_posedge       	: std_ulogic := '0';
        variable Tviol_TMDSch2p_TMDSclkp_negedge 	: std_ulogic := '0';
        variable Tviol_TMDSch2n_TMDSclkp_posedge     	: std_ulogic := '0';
        variable Tviol_TMDSch2n_TMDSclkp_negedge        : std_ulogic := '0';

        variable Tmkr_TMDSch0p_TMDSclkp_posedge        	: VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_TMDSch0p_TMDSclkp_negedge 	: VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_TMDSch0n_TMDSclkp_posedge		: VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_TMDSch0n_TMDSclkp_negedge	        : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_TMDSch1p_TMDSclkp_posedge        	: VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_TMDSch1p_TMDSclkp_negedge 	: VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_TMDSch1n_TMDSclkp_posedge		: VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_TMDSch1n_TMDSclkp_negedge	        : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_TMDSch2p_TMDSclkp_posedge        	: VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_TMDSch2p_TMDSclkp_negedge 	: VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_TMDSch2n_TMDSclkp_posedge		: VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_TMDSch2n_TMDSclkp_negedge	        : VitalTimingDataType := VitalTimingDataInit;

 begin
    if (TimingChecksOn) then

        VitalSetupHoldCheck (
        Violation      => Tviol_TMDSch0p_TMDSclkp_posedge,
        TimingData     => Tmkr_TMDSch0p_TMDSclkp_posedge,
        TestSignal     => TMDSch0p_ipd,
        TestSignalName => "TMDSch0p",
        RefSignal      => TMDSclkp_ipd,
        RefSignalName  => "TMDSclkp",
        SetupHigh      => tsetup_TMDSch0p_TMDSclkp_posedge_posedge,
        SetupLow       => tsetup_TMDSch0p_TMDSclkp_negedge_posedge,
        HoldLow        => thold_TMDSch0p_TMDSclkp_posedge_posedge, 
        HoldHigh       => thold_TMDSch0p_TMDSclkp_negedge_posedge, 
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_TMDS_Deserializer",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);


        VitalSetupHoldCheck (
        Violation      => Tviol_TMDSch0p_TMDSclkp_negedge,
        TimingData     => Tmkr_TMDSch0p_TMDSclkp_negedge,
        TestSignal     => TMDSch0p_ipd,
        TestSignalName => "TMDSch0p",
        RefSignal      => TMDSclkp_ipd,
        RefSignalName  => "TMDSclkp",
        SetupHigh      => tsetup_TMDSch0p_TMDSclkp_posedge_negedge,
        SetupLow       => tsetup_TMDSch0p_TMDSclkp_negedge_negedge,
        HoldLow        => thold_TMDSch0p_TMDSclkp_posedge_negedge, 
        HoldHigh       => thold_TMDSch0p_TMDSclkp_negedge_negedge, 
        CheckEnabled   => true,
        RefTransition  => 'F',
        HeaderMsg      => "/SB_TMDS_Deserializer",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);


        VitalSetupHoldCheck (
        Violation      => Tviol_TMDSch0n_TMDSclkp_posedge,
        TimingData     => Tmkr_TMDSch0n_TMDSclkp_posedge,
        TestSignal     => TMDSch0n_ipd,
        TestSignalName => "TMDSch0n",
        RefSignal      => TMDSclkp_ipd,
        RefSignalName  => "TMDSclkp",
        SetupHigh      => tsetup_TMDSch0n_TMDSclkp_posedge_posedge,
        SetupLow       => tsetup_TMDSch0n_TMDSclkp_negedge_posedge,
        HoldLow        => thold_TMDSch0n_TMDSclkp_posedge_posedge, 
        HoldHigh       => thold_TMDSch0n_TMDSclkp_negedge_posedge, 
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_TMDS_Deserializer",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);


        VitalSetupHoldCheck (
        Violation      => Tviol_TMDSch0n_TMDSclkp_negedge,
        TimingData     => Tmkr_TMDSch0n_TMDSclkp_negedge,
        TestSignal     => TMDSch0n_ipd,
        TestSignalName => "TMDSch0n",
        RefSignal      => TMDSclkp_ipd,
        RefSignalName  => "TMDSclkp",
        SetupHigh      => tsetup_TMDSch0n_TMDSclkp_posedge_negedge,
        SetupLow       => tsetup_TMDSch0n_TMDSclkp_negedge_negedge,
        HoldLow        => thold_TMDSch0n_TMDSclkp_posedge_negedge, 
        HoldHigh       => thold_TMDSch0n_TMDSclkp_negedge_negedge, 
        CheckEnabled   => true,
        RefTransition  => 'F',
        HeaderMsg      => "/SB_TMDS_Deserializer",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);


        VitalSetupHoldCheck (
        Violation      => Tviol_TMDSch1p_TMDSclkp_posedge,
        TimingData     => Tmkr_TMDSch1p_TMDSclkp_posedge,
        TestSignal     => TMDSch1p_ipd,
        TestSignalName => "TMDSch1p",
        RefSignal      => TMDSclkp_ipd,
        RefSignalName  => "TMDSclkp",
        SetupHigh      => tsetup_TMDSch1p_TMDSclkp_posedge_posedge,
        SetupLow       => tsetup_TMDSch1p_TMDSclkp_negedge_posedge,
        HoldLow        => thold_TMDSch1p_TMDSclkp_posedge_posedge, 
        HoldHigh       => thold_TMDSch1p_TMDSclkp_negedge_posedge, 
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_TMDS_Deserializer",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);


        VitalSetupHoldCheck (
        Violation      => Tviol_TMDSch1p_TMDSclkp_negedge,
        TimingData     => Tmkr_TMDSch1p_TMDSclkp_negedge,
        TestSignal     => TMDSch1p_ipd,
        TestSignalName => "TMDSch1p",
        RefSignal      => TMDSclkp_ipd,
        RefSignalName  => "TMDSclkp",
        SetupHigh      => tsetup_TMDSch1p_TMDSclkp_posedge_negedge,
        SetupLow       => tsetup_TMDSch1p_TMDSclkp_negedge_negedge,
        HoldLow        => thold_TMDSch1p_TMDSclkp_posedge_negedge, 
        HoldHigh       => thold_TMDSch1p_TMDSclkp_negedge_negedge, 
        CheckEnabled   => true,
        RefTransition  => 'F',
        HeaderMsg      => "/SB_TMDS_Deserializer",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);


        VitalSetupHoldCheck (
        Violation      => Tviol_TMDSch1n_TMDSclkp_posedge,
        TimingData     => Tmkr_TMDSch1n_TMDSclkp_posedge,
        TestSignal     => TMDSch1n_ipd,
        TestSignalName => "TMDSch1n",
        RefSignal      => TMDSclkp_ipd,
        RefSignalName  => "TMDSclkp",
        SetupHigh      => tsetup_TMDSch1n_TMDSclkp_posedge_posedge,
        SetupLow       => tsetup_TMDSch1n_TMDSclkp_negedge_posedge,
        HoldLow        => thold_TMDSch1n_TMDSclkp_posedge_posedge, 
        HoldHigh       => thold_TMDSch1n_TMDSclkp_negedge_posedge, 
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_TMDS_Deserializer",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);


        VitalSetupHoldCheck (
        Violation      => Tviol_TMDSch1n_TMDSclkp_negedge,
        TimingData     => Tmkr_TMDSch1n_TMDSclkp_negedge,
        TestSignal     => TMDSch1n_ipd,
        TestSignalName => "TMDSch1n",
        RefSignal      => TMDSclkp_ipd,
        RefSignalName  => "TMDSclkp",
        SetupHigh      => tsetup_TMDSch1n_TMDSclkp_posedge_negedge,
        SetupLow       => tsetup_TMDSch1n_TMDSclkp_negedge_negedge,
        HoldLow        => thold_TMDSch1n_TMDSclkp_posedge_negedge, 
        HoldHigh       => thold_TMDSch1n_TMDSclkp_negedge_negedge, 
        CheckEnabled   => true,
        RefTransition  => 'F',
        HeaderMsg      => "/SB_TMDS_Deserializer",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);

        VitalSetupHoldCheck (
        Violation      => Tviol_TMDSch2p_TMDSclkp_posedge,
        TimingData     => Tmkr_TMDSch2p_TMDSclkp_posedge,
        TestSignal     => TMDSch2p_ipd,
        TestSignalName => "TMDSch2p",
        RefSignal      => TMDSclkp_ipd,
        RefSignalName  => "TMDSclkp",
        SetupHigh      => tsetup_TMDSch2p_TMDSclkp_posedge_posedge,
        SetupLow       => tsetup_TMDSch2p_TMDSclkp_negedge_posedge,
        HoldLow        => thold_TMDSch2p_TMDSclkp_posedge_posedge, 
        HoldHigh       => thold_TMDSch2p_TMDSclkp_negedge_posedge, 
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_TMDS_Deserializer",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);


        VitalSetupHoldCheck (
        Violation      => Tviol_TMDSch2p_TMDSclkp_negedge,
        TimingData     => Tmkr_TMDSch2p_TMDSclkp_negedge,
        TestSignal     => TMDSch2p_ipd,
        TestSignalName => "TMDSch2p",
        RefSignal      => TMDSclkp_ipd,
        RefSignalName  => "TMDSclkp",
        SetupHigh      => tsetup_TMDSch2p_TMDSclkp_posedge_negedge,
        SetupLow       => tsetup_TMDSch2p_TMDSclkp_negedge_negedge,
        HoldLow        => thold_TMDSch2p_TMDSclkp_posedge_negedge, 
        HoldHigh       => thold_TMDSch2p_TMDSclkp_negedge_negedge, 
        CheckEnabled   => true,
        RefTransition  => 'F',
        HeaderMsg      => "/SB_TMDS_Deserializer",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);


        VitalSetupHoldCheck (
        Violation      => Tviol_TMDSch2n_TMDSclkp_posedge,
        TimingData     => Tmkr_TMDSch2n_TMDSclkp_posedge,
        TestSignal     => TMDSch2n_ipd,
        TestSignalName => "TMDSch2n",
        RefSignal      => TMDSclkp_ipd,
        RefSignalName  => "TMDSclkp",
        SetupHigh      => tsetup_TMDSch2n_TMDSclkp_posedge_posedge,
        SetupLow       => tsetup_TMDSch2n_TMDSclkp_negedge_posedge,
        HoldLow        => thold_TMDSch2n_TMDSclkp_posedge_posedge, 
        HoldHigh       => thold_TMDSch2n_TMDSclkp_negedge_posedge, 
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_TMDS_Deserializer",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);


        VitalSetupHoldCheck (
        Violation      => Tviol_TMDSch2n_TMDSclkp_negedge,
        TimingData     => Tmkr_TMDSch2n_TMDSclkp_negedge,
        TestSignal     => TMDSch2n_ipd,
        TestSignalName => "TMDSch2n",
        RefSignal      => TMDSclkp_ipd,
        RefSignalName  => "TMDSclkp",
        SetupHigh      => tsetup_TMDSch2n_TMDSclkp_posedge_negedge,
        SetupLow       => tsetup_TMDSch2n_TMDSclkp_negedge_negedge,
        HoldLow        => thold_TMDSch2n_TMDSclkp_posedge_negedge, 
        HoldHigh       => thold_TMDSch2n_TMDSclkp_negedge_negedge, 
        CheckEnabled   => true,
        RefTransition  => 'F',
        HeaderMsg      => "/SB_TMDS_Deserializer",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);
 end if;
end process VITALTimingCheck;


-----------------------------------------------------------------
--VITAL Path Delay
------------------------------------------------------------------
       VITALPathDelay  : process (RAWDATAch0_zd, RAWDATAch1_zd, RAWDATAch2_zd , PLLOUTGLOBALclkx1_zd, PLLOUTCOREclkx1_zd, PLLOUTGLOBALclkx5_zd, PLLOUTCOREclkx5_zd, PLLlock_zd, SDO_zd )

        variable RAWDATAch0_0_GlitchData : VitalGlitchDataType;
        variable RAWDATAch0_1_GlitchData : VitalGlitchDataType;
        variable RAWDATAch0_2_GlitchData : VitalGlitchDataType;
        variable RAWDATAch0_3_GlitchData : VitalGlitchDataType;
        variable RAWDATAch0_4_GlitchData : VitalGlitchDataType;
        variable RAWDATAch0_5_GlitchData : VitalGlitchDataType;
        variable RAWDATAch0_6_GlitchData : VitalGlitchDataType;
        variable RAWDATAch0_7_GlitchData : VitalGlitchDataType;
        variable RAWDATAch0_8_GlitchData : VitalGlitchDataType;
        variable RAWDATAch0_9_GlitchData : VitalGlitchDataType;
        variable RAWDATAch1_0_GlitchData : VitalGlitchDataType;
        variable RAWDATAch1_1_GlitchData : VitalGlitchDataType;
        variable RAWDATAch1_2_GlitchData : VitalGlitchDataType;
        variable RAWDATAch1_3_GlitchData : VitalGlitchDataType;
        variable RAWDATAch1_4_GlitchData : VitalGlitchDataType;
        variable RAWDATAch1_5_GlitchData : VitalGlitchDataType;
        variable RAWDATAch1_6_GlitchData : VitalGlitchDataType;
        variable RAWDATAch1_7_GlitchData : VitalGlitchDataType;
        variable RAWDATAch1_8_GlitchData : VitalGlitchDataType;
        variable RAWDATAch1_9_GlitchData : VitalGlitchDataType;
        variable RAWDATAch2_0_GlitchData : VitalGlitchDataType;
        variable RAWDATAch2_1_GlitchData : VitalGlitchDataType;
        variable RAWDATAch2_2_GlitchData : VitalGlitchDataType;
        variable RAWDATAch2_3_GlitchData : VitalGlitchDataType;
        variable RAWDATAch2_4_GlitchData : VitalGlitchDataType;
        variable RAWDATAch2_5_GlitchData : VitalGlitchDataType;
        variable RAWDATAch2_6_GlitchData : VitalGlitchDataType;
        variable RAWDATAch2_7_GlitchData : VitalGlitchDataType;
        variable RAWDATAch2_8_GlitchData : VitalGlitchDataType;
        variable RAWDATAch2_9_GlitchData : VitalGlitchDataType;

        variable PLLOUTGLOBALclkx1_GlitchData : VitalGlitchDataType;
        variable PLLOUTCOREclkx1_GlitchData : VitalGlitchDataType;
        variable PLLOUTGLOBALclkx5_GlitchData : VitalGlitchDataType;
	variable PLLOUTCOREclkx5_GlitchData: VitalGlitchDataType;
	variable PLLlock_GlitchData : VitalGlitchDataType;
	variable SDO_GlitchData : VitalGlitchDataType;

  begin

      VitalPathDelay01 (
      OutSignal                 => RAWDATAch0(0),
      GlitchData                => RAWDATAch0_0_GlitchData,
      OutSignalName             => "RAWDATAch0(0)",
      OutTemp                   => RAWDATAch0_zd(0),
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_RAWDATAch0_posedge(0),true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => RAWDATAch0(1),
      GlitchData                => RAWDATAch0_1_GlitchData,
      OutSignalName             => "RAWDATAch0(1)",
      OutTemp                   => RAWDATAch0_zd(1),
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_RAWDATAch0_posedge(1),true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => RAWDATAch0(2),
      GlitchData                => RAWDATAch0_2_GlitchData,
      OutSignalName             => "RAWDATAch0(2)",
      OutTemp                   => RAWDATAch0_zd(2),
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_RAWDATAch0_posedge(2),true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => RAWDATAch0(3),
      GlitchData                => RAWDATAch0_3_GlitchData,
      OutSignalName             => "RAWDATAch0(3)",
      OutTemp                   => RAWDATAch0_zd(3),
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_RAWDATAch0_posedge(3),true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => RAWDATAch0(4),
      GlitchData                => RAWDATAch0_4_GlitchData,
      OutSignalName             => "RAWDATAch0(4)",
      OutTemp                   => RAWDATAch0_zd(4),
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_RAWDATAch0_posedge(4),true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => RAWDATAch0(5),
      GlitchData                => RAWDATAch0_5_GlitchData,
      OutSignalName             => "RAWDATAch0(5)",
      OutTemp                   => RAWDATAch0_zd(5),
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_RAWDATAch0_posedge(5),true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => RAWDATAch0(6),
      GlitchData                => RAWDATAch0_6_GlitchData,
      OutSignalName             => "RAWDATAch0(6)",
      OutTemp                   => RAWDATAch0_zd(6),
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_RAWDATAch0_posedge(6),true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => RAWDATAch0(7),
      GlitchData                => RAWDATAch0_7_GlitchData,
      OutSignalName             => "RAWDATAch0(7)",
      OutTemp                   => RAWDATAch0_zd(7),
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_RAWDATAch0_posedge(7),true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => RAWDATAch0(8),
      GlitchData                => RAWDATAch0_8_GlitchData,
      OutSignalName             => "RAWDATAch0(8)",
      OutTemp                   => RAWDATAch0_zd(8),
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_RAWDATAch0_posedge(8),true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => RAWDATAch0(9),
      GlitchData                => RAWDATAch0_9_GlitchData,
      OutSignalName             => "RAWDATAch0(9)",
      OutTemp                   => RAWDATAch0_zd(9),
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_RAWDATAch0_posedge(9),true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => RAWDATAch1(0),
      GlitchData                => RAWDATAch1_0_GlitchData,
      OutSignalName             => "RAWDATAch1(0)",
      OutTemp                   => RAWDATAch1_zd(0),
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_RAWDATAch1_posedge(0),true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => RAWDATAch1(1),
      GlitchData                => RAWDATAch1_1_GlitchData,
      OutSignalName             => "RAWDATAch1(1)",
      OutTemp                   => RAWDATAch1_zd(1),
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_RAWDATAch1_posedge(1),true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => RAWDATAch1(2),
      GlitchData                => RAWDATAch1_2_GlitchData,
      OutSignalName             => "RAWDATAch1(2)",
      OutTemp                   => RAWDATAch1_zd(2),
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_RAWDATAch1_posedge(2),true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => RAWDATAch1(3),
      GlitchData                => RAWDATAch1_3_GlitchData,
      OutSignalName             => "RAWDATAch1(3)",
      OutTemp                   => RAWDATAch1_zd(3),
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_RAWDATAch1_posedge(3),true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => RAWDATAch1(4),
      GlitchData                => RAWDATAch1_4_GlitchData,
      OutSignalName             => "RAWDATAch1(4)",
      OutTemp                   => RAWDATAch1_zd(4),
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_RAWDATAch1_posedge(4),true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => RAWDATAch1(5),
      GlitchData                => RAWDATAch1_5_GlitchData,
      OutSignalName             => "RAWDATAch1(5)",
      OutTemp                   => RAWDATAch1_zd(5),
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_RAWDATAch1_posedge(5),true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => RAWDATAch1(6),
      GlitchData                => RAWDATAch1_6_GlitchData,
      OutSignalName             => "RAWDATAch1(6)",
      OutTemp                   => RAWDATAch1_zd(6),
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_RAWDATAch1_posedge(6),true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => RAWDATAch1(7),
      GlitchData                => RAWDATAch1_7_GlitchData,
      OutSignalName             => "RAWDATAch1(7)",
      OutTemp                   => RAWDATAch1_zd(7),
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_RAWDATAch1_posedge(7),true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => RAWDATAch1(8),
      GlitchData                => RAWDATAch1_8_GlitchData,
      OutSignalName             => "RAWDATAch1(8)",
      OutTemp                   => RAWDATAch1_zd(8),
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_RAWDATAch1_posedge(8),true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => RAWDATAch1(9),
      GlitchData                => RAWDATAch1_9_GlitchData,
      OutSignalName             => "RAWDATAch1(9)",
      OutTemp                   => RAWDATAch1_zd(9),
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_RAWDATAch1_posedge(9),true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => RAWDATAch2(0),
      GlitchData                => RAWDATAch2_0_GlitchData,
      OutSignalName             => "RAWDATAch2(0)",
      OutTemp                   => RAWDATAch2_zd(0),
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_RAWDATAch2_posedge(0),true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => RAWDATAch2(1),
      GlitchData                => RAWDATAch2_1_GlitchData,
      OutSignalName             => "RAWDATAch2(1)",
      OutTemp                   => RAWDATAch2_zd(1),
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_RAWDATAch2_posedge(1),true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => RAWDATAch2(2),
      GlitchData                => RAWDATAch2_2_GlitchData,
      OutSignalName             => "RAWDATAch2(2)",
      OutTemp                   => RAWDATAch2_zd(2),
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_RAWDATAch2_posedge(2),true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => RAWDATAch2(3),
      GlitchData                => RAWDATAch2_3_GlitchData,
      OutSignalName             => "RAWDATAch2(3)",
      OutTemp                   => RAWDATAch2_zd(3),
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_RAWDATAch2_posedge(3),true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => RAWDATAch2(4),
      GlitchData                => RAWDATAch2_4_GlitchData,
      OutSignalName             => "RAWDATAch2(4)",
      OutTemp                   => RAWDATAch2_zd(4),
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_RAWDATAch2_posedge(4),true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => RAWDATAch2(5),
      GlitchData                => RAWDATAch2_5_GlitchData,
      OutSignalName             => "RAWDATAch2(5)",
      OutTemp                   => RAWDATAch2_zd(5),
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_RAWDATAch2_posedge(5),true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => RAWDATAch2(6),
      GlitchData                => RAWDATAch2_6_GlitchData,
      OutSignalName             => "RAWDATAch2(6)",
      OutTemp                   => RAWDATAch2_zd(6),
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_RAWDATAch2_posedge(6),true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => RAWDATAch2(7),
      GlitchData                => RAWDATAch2_7_GlitchData,
      OutSignalName             => "RAWDATAch2(7)",
      OutTemp                   => RAWDATAch2_zd(7),
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_RAWDATAch2_posedge(7),true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => RAWDATAch2(8),
      GlitchData                => RAWDATAch2_8_GlitchData,
      OutSignalName             => "RAWDATAch2(8)",
      OutTemp                   => RAWDATAch2_zd(8),
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_RAWDATAch2_posedge(8),true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => RAWDATAch2(9),
      GlitchData                => RAWDATAch2_9_GlitchData,
      OutSignalName             => "RAWDATAch2(9)",
      OutTemp                   => RAWDATAch2_zd(9),
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_RAWDATAch2_posedge(9),true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => PLLOUTGLOBALclkx1,
      GlitchData                => PLLOUTGLOBALclkx1_GlitchData,
      OutSignalName             => "PLLOUTGLOBALclkx1",
      OutTemp                   => PLLOUTGLOBALclkx1_zd,
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_PLLOUTGLOBALclkx1, true)
                                   ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);


      VitalPathDelay01 (
      OutSignal                 => PLLOUTCOREclkx1,
      GlitchData                => PLLOUTCOREclkx1_GlitchData,
      OutSignalName             => "PLLOUTCOREclkx1",
      OutTemp                   => PLLOUTCOREclkx1_zd,
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_PLLOUTCOREclkx1, true)
                                   ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);


      VitalPathDelay01 (
      OutSignal                 => PLLOUTGLOBALclkx5,
      GlitchData                => PLLOUTGLOBALclkx5_GlitchData,
      OutSignalName             => "PLLOUTGLOBALclkx5",
      OutTemp                   => PLLOUTGLOBALclkx5_zd,
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event, tpd_TMDSclkp_PLLOUTGLOBALclkx5, true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);


      VitalPathDelay01 (
      OutSignal                 => PLLOUTCOREclkx5,
      GlitchData                => PLLOUTCOREclkx5_GlitchData,
      OutSignalName             => "PLLOUTCOREclkx5",
      OutTemp                   => PLLOUTCOREclkx5_zd,
      Paths                     => ( 0 => (TMDSclkp_ipd'last_event,tpd_TMDSclkp_PLLOUTCOREclkx5 , true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

end process VITALPathDelay;

end SB_TMDS_deserializer_V; 

--------------------------------------------------- 
--- 		dvi_deserializer 		 --
---------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;	 
library work;
use work.std_logic_SBT.all;	   

entity dvi_deserializer is
	port ( 
		en  	: in 	std_logic ; 							
		rstn  	: in 	std_logic ; 
		din		: in	std_logic ; 
		clkx5in	: in	std_logic ; 	
		clkx1in	: in 	std_logic ; 
		rawdata : out  	std_logic_vector(9 downto 0)	
	   	  ); 	
end dvi_deserializer;  

architecture dvi_deserializer_arch of dvi_deserializer is	

component mem4x10 is 
	port (
  			WDATAIN	 	: in  	std_logic_vector( 9 downto 0); 
  			WCLK 		: in	std_logic ; 
  			WE		 	: in	std_logic ; 
  			WADDR	 	: in	std_logic_vector(1 downto 0) ; 
  			RADDR	 	: in	std_logic_vector(1 downto 0) ; 
  		    	RDATAOUT 	: out 	std_logic_vector(9 downto 0)
		); 
end component; 		

	type StateType is (ST0,ST1,ST2,ST3,ST4);
    	signal 	n_state ,p_state : StateType;  
  
	
	signal clkx1 , clkx5  		: 	std_logic ; 
	signal din_n0, din_n1  		: 	std_logic ;
	signal 	din_p0			: 	std_logic ; 
	signal 	datain			: 	std_logic_vector( 9 downto 0) ; 
	signal  datain_q		: 	std_logic_vector( 9 downto 0) ;
	signal  mem_rdout		: 	std_logic_vector( 9 downto 0) ;	
	
	signal  pulse_5cnt		: 	std_logic ;
 	signal  sync_wren		: 	std_logic ;
	 
	signal sync_rden		: 	std_logic_vector(3 downto 0);  
	signal rstsync_w		: 	std_logic;  
	signal rstsync_r 		: 	std_logic ;  
	signal wa_rst , ra_rst		: 	std_logic ;						
	
	signal wa			: 	std_logic_vector(1 downto 0) ; 
  	signal ra			: 	std_logic_vector(1 downto 0) ; 

begin

	clkx1 <= ( clkx1in and en ) ; 
	clkx5 <= ( clkx5in and en ) ; 
------------ Data Sampling Section  --------------- 
 	din_n0_proc : process(clkx5,en) 
 	begin 	    
		  if falling_edge(clkx5) then 
			  if(en = '1') then 
				  din_n0 <= din;
		  end if; 
	  end if ; 		  
 	end process din_n0_proc; 	

	din_n1_proc : process(clkx5) 
	begin 
		if rising_edge(clkx5) then 
			din_n1    <= not(din_n0);	
			datain(8) <= din_n1; 
			datain(6) <= datain(8); 
			datain(4) <= datain(6); 
			datain(2) <= datain(4); 
			datain(0) <= datain(2); 
		end  if; 
	end process  din_n1_proc; 

	--always@(posedge clkx5) 
	din_p0_proc : process(clkx5) 
	begin 
		if rising_edge(clkx5) then 
			din_p0 <= din; 
			datain(9) <= not(din_p0); 
			datain(7) <= datain(9); 	
			datain(5) <= datain(7); 
			datain(3) <= datain(5); 
			datain(1) <= datain(3); 
	 	end if; 
	end process  din_p0_proc; 


	datainq_proc : process(clkx5) 
	begin 
		if rising_edge(clkx5) then 
			datain_q<=datain; 		
	 	end if; 
	end process  datainq_proc; 


 	-- State Machine ---- 			  
  statemach_comb: process(p_state,rstn) 
  begin 
	  case p_state  is 
		  when ST0 => 
		  			if (rstn ='1') then 
			  			n_state <= ST1;
		  			else 
						 n_state <= ST0;
		  			end if;  
		  when ST1 => 
		  			if (rstn = '1') then  
						  n_state <= ST2;
					else 
						  n_state <= ST1;
		  			end if;  	   
		  
		  when ST2 => 
		  			if (rstn = '1') then  
						 n_state <= ST3;
					else 
						 n_state <= ST2;
		  			end if;  
		  when ST3 => 
		  			if (rstn = '1') then 
		  				n_state <= ST4; 
					else 
						 n_state <= ST3;
		  			end if;  
		  when others =>  n_state <=ST0; 
	  end case; 
  end process statemach_comb ; 
  
  statemach_seq : process( clkx5,rstn,en ) 
  begin 
	  if(rstn = '0') then
		  	 p_state <= ST0; 
	  elsif  rising_edge(clkx5) then 
		  if (en ='1') then 
			  p_state <= n_state; 
		  end if; 
	  end if; 
 end process statemach_seq; 
 
  with p_state select  
 		pulse_5cnt <= '1' when ST3,
 					  '0' when others; 	 

	 	
 process(clkx5) 
 begin 
	if rising_edge(clkx5) then 
	 sync_wren <= pulse_5cnt;  
	end if; 
 end process; 
 				   
  -- syncronous read , write reset signal gen 
  
  sync_wrrst_proc : process(clkx5)
  begin 									  
	if rising_edge(clkx5)  then 
	  rstsync_w <= rstn; 
	  rstsync_r <= rstsync_w; 
	  wa_rst    <= rstsync_r;	
	  end if ; 
  end process sync_wrrst_proc; 					   
  
   --  delay ra_rst 
  sync_rdrst_proc : process(clkx5)
  begin 									  
	if rising_edge(clkx5)  then    
		sync_rden(0) <= rstsync_r;   
  		sync_rden(1) <= sync_rden(0);
		sync_rden(2) <= sync_rden(1);
		sync_rden(3) <= sync_rden(2);
		ra_rst <= sync_rden(3); 
  	end if ;
  end process sync_rdrst_proc;   
  
  --Address Generation Logics   
  
  wagen_proc : process ( clkx5, wa_rst) 
  begin 
	 if(wa_rst = '0') 	then 	
		  wa <= (others => '0') ; 
	 elsif  rising_edge (clkx5) then 
		 if (sync_wren = '1') then 
			wa <= wa +1 ;  
		 end if; 
	 end if;  
	
  end process wagen_proc; 
		
  rdgen_proc : process (clkx1, ra_rst) 
  begin 								   
	  if(ra_rst = '0') then  
		  ra <= (others => '0') ;  
	  elsif rising_edge(clkx1) then 
  	 	ra <= ra +1;  
	  end if ; 	   
  end process rdgen_proc;  	    
  
  mem4x10_i  : mem4x10   port map (
  			WDATAIN	 => datain_q,
  			WCLK 	 => clkx5,
  			WE	 => sync_wren,
  			WADDR	 => wa,
  			RADDR	 => ra, 
  		    	RDATAOUT => mem_rdout
  								); 
  

 process(clkx1)						  
 begin
	 if rising_edge(clkx1) then 
    		rawdata<=mem_rdout;
	 end if ; 	
 end process; 		  

end dvi_deserializer_arch;

------------------------------------------
----	 clkdelay16  		     -----
------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;	 
library work;
use work.std_logic_SBT.all;	   

entity clkdelay16 is 
	generic (
			BUF_DELAY : time  		:= 100 ps  
		); 		
	port    ( 
			dlyin    : in 	 	std_logic;  
			dlyout	 : out 		std_logic ;  
			dly_sel	 : in 		std_logic_vector( 3 downto 0)
		); 															  	
end clkdelay16;

			
architecture clkdelay16_arch of clkdelay16 is
	signal buf_y   : std_logic_vector( 15 downto 0); 
	signal delayed_data : std_logic; 
begin
 	buf_y(0)  <= dlyin; 
  
	delaytap_gen: for N in 1 to 15 generate
        	buf_y(N) <= buf_y(N-1) after  BUF_DELAY ;             -- 100ps +-25ps.
      	end generate;

      	seldelay_proc: process(dly_sel,buf_y )
        begin
                delayed_data <=buf_y(slv_to_integer(dly_sel));
        end process;

        dlyout <= delayed_data;	 

end clkdelay16_arch;

------------------------------------
----       mem4x10               ---
------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;	 
library work;
use work.std_logic_SBT.all;	   

entity mem4x10  is 
	port 
	(
	WDATAIN 	: in 	std_logic_vector(9 downto 0) ; 
	WCLK		: in	std_logic ; 
	WE			: in	std_logic ; 
	WADDR		: in	std_logic_vector(1 downto 0) ;
	RADDR		: in	std_logic_vector(1 downto 0) ; 
	RDATAOUT	: out 	std_logic_vector(9 downto 0) 
	); 
	
end mem4x10; 

architecture mem4x10_arch of mem4x10 is 

	type ramtype is array (0 to 3) of std_logic_vector (9 downto 0); 
	signal mem : ramtype ; 
	
begin 	
	
	-- read first memory 
	ramwr_proc : process(WCLK) 
   	begin 		
		if rising_edge(WCLK) then 
			if (WE ='1') then 
			mem(conv_integer(unsigned(WADDR))) <= WDATAIN; 								
			end if; 
		end if; 	
    	end process ramwr_proc; 	
	
	RDATAOUT <= mem(conv_integer(unsigned(RADDR))) ;     	
	
end mem4x10_arch;  

----------------------------------------------------------------------------
----			SB_MIPI_RX_2LANE				---- 
----------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;

entity  SB_MIPI_RX_2LANE is 
	generic  (
	
		----------------------------------------------------------------------------------
	        --VITAL PARAMETER
		---------------------------------------------------------------------------------
        	TimingChecksOn  	: boolean := true;
        	Xon   			: boolean := true;
    		MsgOn 			: boolean := false;
        	--- VITAL input port delay 
        	tipd_ENPDESER	  			: VitalDelayType01 := (0 ns, 0 ns);
        	tipd_PU        				: VitalDelayType01 := (0 ns, 0 ns);
        	tipd_DP0 	       			: VitalDelayType01 := (0 ns, 0 ns);
        	tipd_DN0 	       			: VitalDelayType01 := (0 ns, 0 ns);
        	tipd_D0TXLPEN 	       			: VitalDelayType01 := (0 ns, 0 ns);
        	tipd_D0DTXLPP 	       			: VitalDelayType01 := (0 ns, 0 ns);
        	tipd_D0DTXLPN 	       			: VitalDelayType01 := (0 ns, 0 ns);
        	tipd_D0RXLPEN 	       			: VitalDelayType01 := (0 ns, 0 ns);
        	tipd_D0CDEN 	       			: VitalDelayType01 := (0 ns, 0 ns);
        	tipd_D0RXHSEN	       			: VitalDelayType01 := (0 ns, 0 ns);
        	tipd_D0HSDESEREN       			: VitalDelayType01 := (0 ns, 0 ns);
        	tipd_DP1 	       			: VitalDelayType01 := (0 ns, 0 ns);
        	tipd_DN1 	       			: VitalDelayType01 := (0 ns, 0 ns);
        	tipd_D1RXLPEN 	       			: VitalDelayType01 := (0 ns, 0 ns);
        	tipd_D1RXHSEN	       			: VitalDelayType01 := (0 ns, 0 ns);
        	tipd_D1HSDESEREN       			: VitalDelayType01 := (0 ns, 0 ns);
        	tipd_CKP 	       			: VitalDelayType01 := (0 ns, 0 ns);
        	tipd_CKN 	       			: VitalDelayType01 := (0 ns, 0 ns);
        	tipd_CLKRXLPEN	       			: VitalDelayType01 := (0 ns, 0 ns);
        	tipd_CLKRXHSEN	       			: VitalDelayType01 := (0 ns, 0 ns);
		-- VITAL Path Delay 	
        	tpd_DP0_D0DRXLPP	           	: VitalDelayType01 := (0 ns, 0 ns);
        	tpd_DN0_D0DRXLPN   	  	     	: VitalDelayType01 := (0 ns, 0 ns);
        	tpd_DP0_D0DCDP		           	: VitalDelayType01 := (0 ns, 0 ns);
        	tpd_DN0_D0DCDN		           	: VitalDelayType01 := (0 ns, 0 ns);
        	tpd_DP1_D1DRXLPP	           	: VitalDelayType01 := (0 ns, 0 ns);
        	tpd_DN1_D1DRXLPN	           	: VitalDelayType01 := (0 ns, 0 ns);
        	tpd_CKP_CLKDRXLPP	           	: VitalDelayType01 := (0 ns, 0 ns);
        	tpd_CKN_CLKDRXLPN	           	: VitalDelayType01 := (0 ns, 0 ns);
		tpd_CKP_CLKHSBYTE			: VitalDelayType01 := (0 ns, 0 ns);
		tpd_CKP_D0HSBYTECLKD			: VitalDelayType01 := (0 ns, 0 ns);	
        	-- VITAL clk-to-output path delay
                tpd_CKP_D0HSRXDATA_posedge 		: VitalDelayArrayType01( 7 downto 0) := (others => (0 ns, 0 ns));
                tpd_CKP_D1HSRXDATA_posedge 		:  VitalDelayArrayType01(7 downto 0) := (others => (0 ns, 0 ns));

		tpd_CKP_D0SYNC_posedge			: VitalDelayType01 := (0 ns, 0 ns);	
		tpd_CKP_D0ERRSYNC_posedge		: VitalDelayType01 := (0 ns, 0 ns);	
		tpd_CKP_D0NOSYNC_negedge		: VitalDelayType01 := (0 ns, 0 ns);	
		tpd_CKP_D1SYNC_posedge			: VitalDelayType01 := (0 ns, 0 ns);	
		tpd_CKP_D1ERRSYNC_posedge		: VitalDelayType01 := (0 ns, 0 ns);	
		tpd_CKP_D1NOSYNC_negedge		: VitalDelayType01 := (0 ns, 0 ns);	

		-- VITAL Setup delays 
	        tsetup_DP0_CKP_posedge_posedge 		: VitalDelayType                   := 0 ns; 
           	tsetup_DP0_CKP_negedge_posedge	 	: VitalDelayType                   := 0 ns; 
	        tsetup_DP0_CKP_posedge_negedge 		: VitalDelayType                   := 0 ns; 
           	tsetup_DP0_CKP_negedge_negedge	 	: VitalDelayType                   := 0 ns; 
	        tsetup_DN0_CKP_posedge_posedge 		: VitalDelayType                   := 0 ns; 
           	tsetup_DN0_CKP_negedge_posedge	 	: VitalDelayType                   := 0 ns; 
	        tsetup_DN0_CKP_posedge_negedge 		: VitalDelayType                   := 0 ns; 
           	tsetup_DN0_CKP_negedge_negedge	 	: VitalDelayType                   := 0 ns; 
	        tsetup_DP1_CKP_posedge_posedge 		: VitalDelayType                   := 0 ns; 
           	tsetup_DP1_CKP_negedge_posedge	 	: VitalDelayType                   := 0 ns; 
	        tsetup_DP1_CKP_posedge_negedge 		: VitalDelayType                   := 0 ns; 
           	tsetup_DP1_CKP_negedge_negedge	 	: VitalDelayType                   := 0 ns; 
	        tsetup_DN1_CKP_posedge_posedge 		: VitalDelayType                   := 0 ns; 
           	tsetup_DN1_CKP_negedge_posedge	 	: VitalDelayType                   := 0 ns; 
	        tsetup_DN1_CKP_posedge_negedge 		: VitalDelayType                   := 0 ns; 
           	tsetup_DN1_CKP_negedge_negedge	 	: VitalDelayType                   := 0 ns; 
		-- VITAL Hold delays 
	        thold_DP0_CKP_posedge_posedge 		: VitalDelayType                   := 0 ns; 
           	thold_DP0_CKP_negedge_posedge	 	: VitalDelayType                   := 0 ns; 
	        thold_DP0_CKP_posedge_negedge 		: VitalDelayType                   := 0 ns; 
           	thold_DP0_CKP_negedge_negedge	 	: VitalDelayType                   := 0 ns; 
	        thold_DN0_CKP_posedge_posedge 		: VitalDelayType                   := 0 ns; 
           	thold_DN0_CKP_negedge_posedge	 	: VitalDelayType                   := 0 ns; 
	        thold_DN0_CKP_posedge_negedge 		: VitalDelayType                   := 0 ns; 
           	thold_DN0_CKP_negedge_negedge	 	: VitalDelayType                   := 0 ns; 
	        thold_DP1_CKP_posedge_posedge 		: VitalDelayType                   := 0 ns; 
           	thold_DP1_CKP_negedge_posedge	 	: VitalDelayType                   := 0 ns; 
	        thold_DP1_CKP_posedge_negedge 		: VitalDelayType                   := 0 ns; 
           	thold_DP1_CKP_negedge_negedge	 	: VitalDelayType                   := 0 ns; 
	        thold_DN1_CKP_posedge_posedge 		: VitalDelayType                   := 0 ns; 
           	thold_DN1_CKP_negedge_posedge	 	: VitalDelayType                   := 0 ns; 
	        thold_DN1_CKP_posedge_negedge 		: VitalDelayType                   := 0 ns; 
           	thold_DN1_CKP_negedge_negedge	 	: VitalDelayType                   := 0 ns 
		); 

	port   ( 
		-- Common Interface Pins 
		ENPDESER	: in 		std_logic ; 	
	  	PU		: in		std_logic ; 
		-- Data0 Interface Pins 
		DP0		: in 		std_logic ; 	
		DN0		: in		std_logic ;
		D0RXHSEN	: in 		std_logic ;
  		D0DTXLPP	: in		std_logic ;
  		D0DTXLPN	: in 		std_logic ;
 		D0TXLPEN 	: in		std_logic ; 
 		D0DRXLPP	: out 		std_logic ; 
  		D0DRXLPN	: out 		std_logic ; 
		D0RXLPEN	: in		std_logic ;
 		D0DCDP		: out		std_logic ;
		D0DCDN		: out 		std_logic ;
		D0CDEN		: in		std_logic ; 
  		D0HSDESEREN 	: in 		std_logic ; 
  		D0HSRXDATA  	: out 		std_logic_vector ( 7 downto 0) ;
	    	D0HSBYTECLKD	: out		std_logic ; 
  		D0SYNC		: out		std_logic ;
  		D0ERRSYNC   	: out		std_logic ;
 		D0NOSYNC	: out		std_logic ;
	 	--  DATA1 Interface Pins
 		DP1 		: in		std_logic ;
 		DN1		: in		std_logic ;
	    	D1RXHSEN	: in		std_logic ;
		D1DRXLPP	: out		std_logic ;
		D1DRXLPN	: out		std_logic ;
	    	D1RXLPEN	: in		std_logic ;
	    	D1HSDESEREN	: in		std_logic ;
 		D1HSRXDATA	: out 		std_logic_vector ( 7 downto 0) ; 
 		D1SYNC		: out 		std_logic ; 
  		D1ERRSYNC	: out 		std_logic ;
  		D1NOSYNC	: out 		std_logic ;
	 	--  CLOCK Interface Pins
 		CKP		: in		std_logic ;
 		CKN		: in		std_logic ;
		CLKRXHSEN	: in		std_logic ;
 		CLKDRXLPP	: out 		std_logic ;
  		CLKDRXLPN	: out 		std_logic ;
 		CLKRXLPEN	: in		std_logic ;
        	CLKHSBYTE 	: out 		std_logic
		); 

	attribute VITAL_LEVEL0 of SB_MIPI_RX_2LANE : entity is true;
	 
end SB_MIPI_RX_2LANE;  

architecture SB_MIPI_RX_2LANE_V of SB_MIPI_RX_2LANE is

  attribute VITAL_LEVEL0 of SB_MIPI_RX_2LANE_V  : architecture is true; 

component X105DSI_RX is 
	 port (
		-- Power &  Common Interface Pins 
	VDDA		: in 		std_logic ; 
	VSSA		: in		std_logic ;
	DVSS		: in		std_logic ;
	ENP_DESER	: in		std_logic ;
	PD		: in 		std_logic ;
	   -- DATA0 Interface pins
	DP0		: inout 	std_logic ;
	DN0		: inout 	std_logic ;
	D0_RXHSEN	: in		std_logic ;
	D0_DTXLPP	: in		std_logic ;
	D0_DTXLPN	: in		std_logic ;
	D0_TXLPEN 	: in		std_logic ;
	D0_DRXLPP	: out		std_logic ;
	D0_DRXLPN	: out 		std_logic ;
	D0_RXLPEN	: in		std_logic ;
	D0_DCDP		: out		std_logic ;
	D0_DCDN		: out		std_logic ;
	D0_CDEN		: in		std_logic ;
	D0_HS_DESER_EN	: in	std_logic ;
	D0_HSRX_DATA	: out	std_logic_vector(7 downto 0) ;
	D0_HS_BYTE_CLKD	: out	std_logic ;
	D0_SYNC		: out 	std_logic ;
	D0_ERRSYNC	: out	std_logic ;
	D0_NOSYNC	: out 	std_logic ;
	   -- DATA1 Lane Interface Pins  
	DP1		: in	std_logic ;
	DN1		: in	std_logic ;
	D1_RXHSEN	: in	std_logic ;
	D1_DRXLPP	: out	std_logic ;
	D1_DRXLPN	: out 	std_logic ;
	D1_RXLPEN	: in	std_logic ;
	D1_HS_DESER_EN	: in	std_logic ;
	D1_HSRX_DATA	: out 	std_logic_vector(7 downto 0) ;
	D1_SYNC		: out 	std_logic ;
	D1_ERRSYNC	: out 	std_logic ;
	D1_NOSYNC	: out	std_logic ;
	
	-- CLOCK Interface Pins
	CKP		: in 	std_logic ;
	CKN		: in    std_logic ;
	CLK_RXHSEN	: in	std_logic ;
	CLK_DRXLPP	: out 	std_logic ;
	CLK_DRXLPN	: out	std_logic ;
	CLK_RXLPEN	: in 	std_logic ;
	CLK_HS_BYTE	: out 	std_logic 
	); 
end component; 

	signal  ENPDESER_ipd	      : std_ulogic := 'X';
        signal  PU_ipd		      : std_ulogic := 'X';
        signal  DP0_ipd               : std_ulogic := 'X';
        signal  DN0_ipd               : std_ulogic := 'X';
        signal  D0TXLPEN_ipd          : std_ulogic := 'X';
        signal  D0DTXLPP_ipd          : std_ulogic := 'X';
        signal  D0DTXLPN_ipd          : std_ulogic := 'X';
        signal  D0RXLPEN_ipd          : std_ulogic := 'X';
        signal  D0CDEN_ipd            : std_ulogic := 'X';
        signal  D0RXHSEN_ipd          : std_ulogic := 'X';
        signal  D0HSDESEREN_ipd       : std_ulogic := 'X';
        signal  DP1_ipd               : std_ulogic := 'X';
        signal  DN1_ipd               : std_ulogic := 'X';
        signal  D1RXLPEN_ipd          : std_ulogic := 'X';
        signal  D1RXHSEN_ipd          : std_ulogic := 'X'; 
        signal  D1HSDESEREN_ipd       : std_ulogic := 'X'; 
        signal  CKP_ipd               : std_ulogic := 'X'; 
        signal  CKN_ipd               : std_ulogic := 'X'; 
        signal  CLKRXLPEN_ipd         : std_ulogic := 'X'; 
        signal  CLKRXHSEN_ipd         : std_ulogic := 'X'; 

	signal	D0DRXLPP_zd	      : std_ulogic ; 
	signal	D0DRXLPN_zd	      : std_ulogic ; 
	signal 	D0DCDP_zd	      : std_ulogic ;
	signal  D0DCDN_zd	      : std_ulogic ; 
	signal  D0HSRXDATA_zd 	      : std_logic_vector( 7 downto 0); 
	signal	D0HSBYTECLKD_zd	      : std_ulogic ;
	signal  D0SYNC_zd	      : std_ulogic ;
	signal  D0ERRSYNC_zd	      : std_ulogic ;
	signal  D0NOSYNC_zd	      : std_ulogic ;

	signal  D1DRXLPP_zd 	      : std_ulogic ;
	signal  D1DRXLPN_zd	      : std_ulogic ;
	signal  D1HSRXDATA_zd	      : std_logic_vector( 7 downto 0);    
	signal  D1SYNC_zd	      : std_ulogic ;
	signal  D1ERRSYNC_zd	      : std_ulogic ;  
	signal  D1NOSYNC_zd	      : std_ulogic ; 

	signal	CLKDRXLPP_zd	      : std_ulogic ;
	signal  CLKDRXLPN_zd	      : std_ulogic ;
	signal  CLKHSBYTE_zd	      : std_ulogic ; 

 
	signal not_PU : std_logic ; 	
	signal in_DP0 : std_logic ;
	signal in_DN0 : std_logic ;  
	signal in_DP1 : std_logic ;
	signal in_DN1 : std_logic ;  
	signal in_CKP : std_logic ;
	signal in_CKN : std_logic ;  
	

begin 

 WireDelay   : block
 begin
          VitalWireDelay (ENPDESER_ipd,ENPDESER, tipd_ENPDESER );
          VitalWireDelay (PU_ipd , PU, tipd_PU );
	  VitalWireDelay (DP0_ipd, DP0, tipd_DP0 ); 
	  VitalWireDelay (DN0_ipd, DN0, tipd_DN0 ); 
	  VitalWireDelay (D0TXLPEN_ipd, D0TXLPEN, tipd_D0TXLPEN ); 
	  VitalWireDelay (D0DTXLPP_ipd, D0DTXLPP, tipd_D0DTXLPP  ); 
	  VitalWireDelay (D0DTXLPN_ipd , D0DTXLPN, tipd_D0DTXLPN  ); 
	  VitalWireDelay (D0RXLPEN_ipd, D0RXLPEN, tipd_D0RXLPEN  ); 
	  VitalWireDelay (D0CDEN_ipd , D0CDEN, tipd_D0CDEN  ); 
	  VitalWireDelay (D0RXHSEN_ipd , D0RXHSEN, tipd_D0RXHSEN  ); 
	  VitalWireDelay (D0HSDESEREN_ipd , D0HSDESEREN, tipd_D0HSDESEREN  ); 
	  VitalWireDelay (DP1_ipd, DP1, tipd_DP1  ); 
	  VitalWireDelay (DN1_ipd, DN1, tipd_DN1  ); 
	  VitalWireDelay (D1RXLPEN_ipd, D1RXLPEN, tipd_D1RXLPEN  ); 
	  VitalWireDelay (D1RXHSEN_ipd, D1RXHSEN, tipd_D1RXHSEN  ); 
	  VitalWireDelay (D1HSDESEREN_ipd , D1HSDESEREN, tipd_D1HSDESEREN );  
	  VitalWireDelay (CKP_ipd, CKP, tipd_CKP  ); 
	  VitalWireDelay (CKN_ipd, CKN, tipd_CKN  ); 
	  VitalWireDelay (CLKRXLPEN_ipd , CLKRXLPEN, tipd_CLKRXLPEN  ); 
	  VitalWireDelay (CLKRXHSEN_ipd, CLKRXHSEN, tipd_CLKRXHSEN   ); 
 end block;

 -- Behavioral sections 
	not_PU <= not(PU_ipd); 
	in_DP0 <= DP0_ipd ; 
	in_DN0 <= DN0_ipd ; 
	in_DP1 <= DP1_ipd ; 
	in_DN1 <= DN1_ipd ;
	in_CKP <= CKP_ipd ;  
	in_CKN <= CKN_ipd ; 
	
u_mipi_slave_analog  : X105DSI_RX   

	port map (
		-- Power and Ground Pins
	  VDDA 		=> '1',
	  VSSA 		=> '0', 
	  DVSS  	=> '0',
	 	-- Common Interface pins 
	  ENP_DESER  	=> ENPDESER_ipd,
	  PD         	=> not_pu , 
	 	-- Data0 Interface pins
	  DP0 		=> in_DP0,
	  DN0           => in_DN0,
	  D0_RXHSEN     => D0RXHSEN_ipd,
	  D0_DTXLPP     => D0DTXLPP_ipd,
	  D0_DTXLPN     => D0DTXLPN_ipd,
	  D0_TXLPEN     => D0TXLPEN_ipd,
	  D0_DRXLPP     => D0DRXLPP_zd,
	  D0_DRXLPN     => D0DRXLPN_zd,
	  D0_RXLPEN     => D0RXLPEN_ipd,
	  D0_DCDP       => D0DCDP_zd,
	  D0_DCDN       => D0DCDN_zd,
	  D0_CDEN       => D0CDEN_ipd,
	  D0_HS_DESER_EN => D0HSDESEREN_ipd,
	  D0_HSRX_DATA   => D0HSRXDATA_zd,
	  D0_HS_BYTE_CLKD => D0HSBYTECLKD_zd,
	  D0_SYNC         => D0SYNC_zd,
	  D0_ERRSYNC      => D0ERRSYNC_zd,
	  D0_NOSYNC       => D0NOSYNC_zd,
	 	-- DATA1 Interface pins
	  DP1             => in_DP1,
	  DN1             => in_DN1,
	  D1_RXHSEN       => D1RXHSEN_ipd,
	  D1_DRXLPP       => D1DRXLPP_zd,
	  D1_DRXLPN       => D1DRXLPN_zd,
	  D1_RXLPEN       => D1RXLPEN_ipd,
	  D1_HS_DESER_EN  => D1HSDESEREN_ipd,
	  D1_HSRX_DATA    => D1HSRXDATA_zd,
	  D1_SYNC         => D1SYNC_zd,
	  D1_ERRSYNC      => D1ERRSYNC_zd,
	  D1_NOSYNC       => D1NOSYNC_zd,
	 	--  CLOCK Interface pins
	  CKP             => in_CKP,
	  CKN             => in_CKN,
	  CLK_RXHSEN      => CLKRXHSEN_ipd,
	  CLK_DRXLPP      => CLKDRXLPP_zd,
	  CLK_DRXLPN      => CLKDRXLPN_zd,
	  CLK_RXLPEN      => CLKRXLPEN_ipd,
	  CLK_HS_BYTE     => CLKHSBYTE_zd
	  );

-------------------------------------------------------------------
--VITAL timing check
------------------------------------------------------------------
  VITALTimingCheck : process (CKP_ipd, DP0_ipd, DN0_ipd, DP1_ipd , DN1_ipd)
        variable Tviol_DP0_CKP_posedge          	: std_ulogic := '0';
        variable Tviol_DN0_CKP_posedge 			: std_ulogic := '0';
        variable Tviol_DP1_CKP_posedge 		    	: std_ulogic := '0';
        variable Tviol_DN1_CKP_posedge 		        : std_ulogic := '0';
        variable Tviol_DP0_CKP_negedge           	: std_ulogic := '0';
        variable Tviol_DN0_CKP_negedge 			: std_ulogic := '0';
        variable Tviol_DP1_CKP_negedge 		    	: std_ulogic := '0';
        variable Tviol_DN1_CKP_negedge 		        : std_ulogic := '0';

        variable Tmkr_DP0_CKP_posedge             	: VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_DN0_CKP_posedge    		: VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_DP1_CKP_posedge     		: VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_DN1_CKP_posedge 		        : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_DP0_CKP_negedge             	: VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_DN0_CKP_negedge    		: VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_DP1_CKP_negedge     		: VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_DN1_CKP_negedge 		        : VitalTimingDataType := VitalTimingDataInit;


 begin
    if (TimingChecksOn) then

        VitalSetupHoldCheck (
        Violation      => Tviol_DP0_CKP_posedge,
        TimingData     => Tmkr_DP0_CKP_posedge,
        TestSignal     => DP0_ipd,
        TestSignalName => "DP0",
        RefSignal      => CKP_ipd,
        RefSignalName  => "CKP",
        SetupHigh      => tsetup_DP0_CKP_posedge_posedge,
        SetupLow       => tsetup_DP0_CKP_negedge_posedge,
        HoldLow        => thold_DP0_CKP_negedge_posedge,
        HoldHigh       => thold_DP0_CKP_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MIPI_RX",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);


        VitalSetupHoldCheck (
        Violation      => Tviol_DN0_CKP_posedge,
        TimingData     => Tmkr_DN0_CKP_posedge,
        TestSignal     => DN0_ipd,
        TestSignalName => "DN0",
        RefSignal      => CKP_ipd,
        RefSignalName  => "CKP",
        SetupHigh      => tsetup_DN0_CKP_posedge_posedge,
        SetupLow       => tsetup_DN0_CKP_negedge_posedge,
        HoldLow        => thold_DN0_CKP_negedge_posedge,
        HoldHigh       => thold_DN0_CKP_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MIPI_RX",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);

        VitalSetupHoldCheck (
        Violation      => Tviol_DP1_CKP_posedge,
        TimingData     => Tmkr_DP1_CKP_posedge,
        TestSignal     => DP1_ipd,
        TestSignalName => "DP1",
        RefSignal      => CKP_ipd,
        RefSignalName  => "CKP",
        SetupHigh      => tsetup_DP1_CKP_posedge_posedge,
        SetupLow       => tsetup_DP1_CKP_negedge_posedge,
        HoldLow        => thold_DP1_CKP_negedge_posedge,
        HoldHigh       => thold_DP1_CKP_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MIPI_RX",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);


        VitalSetupHoldCheck (
        Violation      => Tviol_DN1_CKP_posedge,
        TimingData     => Tmkr_DN1_CKP_posedge,
        TestSignal     => DN1_ipd,
        TestSignalName => "DN1",
        RefSignal      => CKP_ipd,
        RefSignalName  => "CKP",
        SetupHigh      => tsetup_DN1_CKP_posedge_posedge,
        SetupLow       => tsetup_DN1_CKP_negedge_posedge,
        HoldLow        => thold_DN1_CKP_negedge_posedge,
        HoldHigh       => thold_DN1_CKP_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MIPI_RX",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);


        VitalSetupHoldCheck (
        Violation      => Tviol_DP0_CKP_negedge,
        TimingData     => Tmkr_DP0_CKP_negedge,
        TestSignal     => DP0_ipd,
        TestSignalName => "DP0",
        RefSignal      => CKP_ipd,
        RefSignalName  => "CKP",
        SetupHigh      => tsetup_DP0_CKP_posedge_negedge,
        SetupLow       => tsetup_DP0_CKP_negedge_negedge,
        HoldLow        => thold_DP0_CKP_negedge_negedge,
        HoldHigh       => thold_DP0_CKP_posedge_negedge,
        CheckEnabled   => true,
        RefTransition  => 'F',
        HeaderMsg      => "/SB_MIPI_RX",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);


        VitalSetupHoldCheck (
        Violation      => Tviol_DN0_CKP_negedge,
        TimingData     => Tmkr_DN0_CKP_negedge,
        TestSignal     => DN0_ipd,
        TestSignalName => "DN0",
        RefSignal      => CKP_ipd,
        RefSignalName  => "CKP",
        SetupHigh      => tsetup_DN0_CKP_posedge_negedge,
        SetupLow       => tsetup_DN0_CKP_negedge_negedge,
        HoldLow        => thold_DN0_CKP_negedge_negedge,
        HoldHigh       => thold_DN0_CKP_posedge_negedge,
        CheckEnabled   => true,
        RefTransition  => 'F',
        HeaderMsg      => "/SB_MIPI_RX",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);

        VitalSetupHoldCheck (
        Violation      => Tviol_DP1_CKP_negedge,
        TimingData     => Tmkr_DP1_CKP_negedge,
        TestSignal     => DP1_ipd,
        TestSignalName => "DP1",
        RefSignal      => CKP_ipd,
        RefSignalName  => "CKP",
        SetupHigh      => tsetup_DP1_CKP_posedge_negedge,
        SetupLow       => tsetup_DP1_CKP_negedge_negedge,
        HoldLow        => thold_DP1_CKP_negedge_negedge,
        HoldHigh       => thold_DP1_CKP_posedge_negedge,
        CheckEnabled   => true,
        RefTransition  => 'F',
        HeaderMsg      => "/SB_MIPI_RX",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);


        VitalSetupHoldCheck (
        Violation      => Tviol_DN1_CKP_negedge,
        TimingData     => Tmkr_DN1_CKP_negedge,
        TestSignal     => DN1_ipd,
        TestSignalName => "DN1",
        RefSignal      => CKP_ipd,
        RefSignalName  => "CKP",
        SetupHigh      => tsetup_DN1_CKP_posedge_negedge,
        SetupLow       => tsetup_DN1_CKP_negedge_negedge,
        HoldLow        => thold_DN1_CKP_negedge_negedge,
        HoldHigh       => thold_DN1_CKP_posedge_negedge,
        CheckEnabled   => true,
        RefTransition  => 'F',
        HeaderMsg      => "/SB_MIPI_RX",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);
 end if;
end process VITALTimingCheck;

-----------------------------------------------------------------
--VITAL Path Delay
------------------------------------------------------------------
       VITALPathDelay  : process (D0DRXLPP_zd,D0DRXLPN_zd,D0DCDP_zd,D0DCDN_zd,D0HSRXDATA_zd, D0HSBYTECLKD_zd,D0SYNC_zd, D0ERRSYNC_zd, D0NOSYNC_zd, D1DRXLPP_zd, D1DRXLPN_zd, D1HSRXDATA_zd, D1SYNC_zd, D1ERRSYNC_zd, D1NOSYNC_zd, CLKDRXLPP_zd, CLKDRXLPN_zd, CLKHSBYTE_zd  )

        variable D0DRXLPP_GlitchData : VitalGlitchDataType;
        variable D0DRXLPN_GlitchData : VitalGlitchDataType;
        variable D0DCDP_GlitchData : VitalGlitchDataType;
        variable D0DCDN_GlitchData : VitalGlitchDataType;
	variable D0HSRXDATA_GlitchData0 : VitalGlitchDataType;
	variable D0HSRXDATA_GlitchData1 : VitalGlitchDataType;
	variable D0HSRXDATA_GlitchData2 : VitalGlitchDataType;
	variable D0HSRXDATA_GlitchData3 : VitalGlitchDataType;
	variable D0HSRXDATA_GlitchData4 : VitalGlitchDataType;
	variable D0HSRXDATA_GlitchData5 : VitalGlitchDataType;
	variable D0HSRXDATA_GlitchData6 : VitalGlitchDataType;
	variable D0HSRXDATA_GlitchData7 : VitalGlitchDataType;
	variable D0HSBYTECLKD_GlitchData : VitalGlitchDataType;
	variable D0SYNC_GlitchData : VitalGlitchDataType;
	variable D0ERRSYNC_GlitchData : VitalGlitchDataType;
	variable D0NOSYNC_GlitchData : VitalGlitchDataType;

	
        variable D1DRXLPP_GlitchData : VitalGlitchDataType;
        variable D1DRXLPN_GlitchData : VitalGlitchDataType;
	variable D1HSRXDATA_GlitchData0 : VitalGlitchDataType;
	variable D1HSRXDATA_GlitchData1 : VitalGlitchDataType;
	variable D1HSRXDATA_GlitchData2 : VitalGlitchDataType;
	variable D1HSRXDATA_GlitchData3 : VitalGlitchDataType;
	variable D1HSRXDATA_GlitchData4 : VitalGlitchDataType;
	variable D1HSRXDATA_GlitchData5 : VitalGlitchDataType;
	variable D1HSRXDATA_GlitchData6 : VitalGlitchDataType;
	variable D1HSRXDATA_GlitchData7 : VitalGlitchDataType;
	variable D1SYNC_GlitchData : VitalGlitchDataType;
	variable D1ERRSYNC_GlitchData : VitalGlitchDataType;
	variable D1NOSYNC_GlitchData : VitalGlitchDataType;

	
	variable CLKDRXLPP_GlitchData : VitalGlitchDataType;
	variable CLKDRXLPN_GlitchData : VitalGlitchDataType;
	variable CLKHSBYTE_GlitchData : VitalGlitchDataType;

  begin

      VitalPathDelay01 (
      OutSignal                 => D0DRXLPP,
      GlitchData                => D0DRXLPP_GlitchData,
      OutSignalName             => "D0DRXLPP",
      OutTemp                   => D0DRXLPP_zd,
      Paths                     => ( 0 => (DP0_ipd'last_event, tpd_DP0_D0DRXLPP, true)
                                   ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);


      VitalPathDelay01 (
      OutSignal                 => D0DRXLPN,
      GlitchData                => D0DRXLPN_GlitchData,
      OutSignalName             => "D0DRXLPN",
      OutTemp                   => D0DRXLPN_zd,
      Paths                     => ( 0 => (DN0_ipd'last_event, tpd_DN0_D0DRXLPN, true)
                                   ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);


      VitalPathDelay01 (
      OutSignal                 => D0DCDP,
      GlitchData                => D0DCDP_GlitchData,
      OutSignalName             => "D0DCDP",
      OutTemp                   => D0DCDP_zd,
      Paths                     => ( 0 => (DP0_ipd'last_event, tpd_DP0_D0DCDP, true)
                                   ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);


      VitalPathDelay01 (
      OutSignal                 => D0DCDN,
      GlitchData                => D0DCDN_GlitchData,
      OutSignalName             => "D0DCDN",
      OutTemp                   => D0DCDN_zd,
      Paths                     => ( 0 => (DN0_ipd'last_event, tpd_DN0_D0DCDN, true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);


      VitalPathDelay01 (
      OutSignal                 => D0HSRXDATA(0),
      GlitchData                => D0HSRXDATA_GlitchData0,
      OutSignalName             => "D0HSRXDATA(0)",
      OutTemp                   => D0HSRXDATA_zd(0),
      Paths                     => ( 0 => (CKP_ipd'last_event,tpd_CKP_D0HSRXDATA_posedge(0) ,true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

	
      VitalPathDelay01 (
      OutSignal                 => D0HSRXDATA(1),
      GlitchData                => D0HSRXDATA_GlitchData1,
      OutSignalName             => "D0HSRXDATA(1)",
      OutTemp                   => D0HSRXDATA_zd(1),
      Paths                     => ( 0 => (CKP_ipd'last_event,tpd_CKP_D0HSRXDATA_posedge(1) ,true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => D0HSRXDATA(2),
      GlitchData                => D0HSRXDATA_GlitchData2,
      OutSignalName             => "D0HSRXDATA(2)",
      OutTemp                   => D0HSRXDATA_zd(2),
      Paths                     => ( 0 => (CKP_ipd'last_event,tpd_CKP_D0HSRXDATA_posedge(2) ,true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => D0HSRXDATA(3),
      GlitchData                => D0HSRXDATA_GlitchData3,
      OutSignalName             => "D0HSRXDATA(3)",
      OutTemp                   => D0HSRXDATA_zd(3),
      Paths                     => ( 0 => (CKP_ipd'last_event,tpd_CKP_D0HSRXDATA_posedge(3) ,true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => D0HSRXDATA(4),
      GlitchData                => D0HSRXDATA_GlitchData4,
      OutSignalName             => "D0HSRXDATA(4)",
      OutTemp                   => D0HSRXDATA_zd(4),
      Paths                     => ( 0 => (CKP_ipd'last_event,tpd_CKP_D0HSRXDATA_posedge(4) ,true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => D0HSRXDATA(5),
      GlitchData                => D0HSRXDATA_GlitchData5,
      OutSignalName             => "D0HSRXDATA(5)",
      OutTemp                   => D0HSRXDATA_zd(5),
      Paths                     => ( 0 => (CKP_ipd'last_event,tpd_CKP_D0HSRXDATA_posedge(5) ,true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => D0HSRXDATA(6),
      GlitchData                => D0HSRXDATA_GlitchData6,
      OutSignalName             => "D0HSRXDATA(6)",
      OutTemp                   => D0HSRXDATA_zd(6),
      Paths                     => ( 0 => (CKP_ipd'last_event,tpd_CKP_D0HSRXDATA_posedge(6) ,true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => D0HSRXDATA(7),
      GlitchData                => D0HSRXDATA_GlitchData7,
      OutSignalName             => "D0HSRXDATA(7)",
      OutTemp                   => D0HSRXDATA_zd(7),
      Paths                     => ( 0 => (CKP_ipd'last_event,tpd_CKP_D0HSRXDATA_posedge(7) ,true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);


      VitalPathDelay01 (
      OutSignal                 => D0HSBYTECLKD,
      GlitchData                => D0HSBYTECLKD_GlitchData,
      OutSignalName             => "D0HSBYTECLKD",
      OutTemp                   => D0HSBYTECLKD_zd,
      Paths                     => ( 0 => (CKP_ipd'last_event, tpd_CKP_D0HSBYTECLKD, true)
                                   ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);


      VitalPathDelay01 (
      OutSignal                 => D0SYNC,
      GlitchData                => D0SYNC_GlitchData,
      OutSignalName             => "D0SYNC",
      OutTemp                   => D0SYNC_zd,
      Paths                     => ( 0 => (CKP_ipd'last_event, tpd_CKP_D0SYNC_posedge, true)),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);


      VitalPathDelay01 (
      OutSignal                 => D0ERRSYNC,
      GlitchData                => D0ERRSYNC_GlitchData,
      OutSignalName             => "D0ERRSYNC",
      OutTemp                   => D0ERRSYNC_zd,
      Paths                     => ( 0 => (CKP_ipd'last_event, tpd_CKP_D0ERRSYNC_posedge, true)),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => D0NOSYNC,
      GlitchData                => D0NOSYNC_GlitchData,
      OutSignalName             => "D0NOSYNC",
      OutTemp                   => D0NOSYNC_zd,
      Paths                     => ( 0 => (CKP_ipd'last_event, tpd_CKP_D0NOSYNC_negedge, true)),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);


      VitalPathDelay01 (
      OutSignal                 => D1DRXLPP,
      GlitchData                => D1DRXLPP_GlitchData,
      OutSignalName             => "D1DRXLPP",
      OutTemp                   => D1DRXLPP_zd,
      Paths                     => ( 0 => (DP1_ipd'last_event, tpd_DP1_D1DRXLPP, true)
                                   ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);


      VitalPathDelay01 (
      OutSignal                 => D1DRXLPN,
      GlitchData                => D1DRXLPN_GlitchData,
      OutSignalName             => "D1DRXLPN",
      OutTemp                   => D1DRXLPN_zd,
      Paths                     => ( 0 => (DN1_ipd'last_event, tpd_DN1_D1DRXLPN, true)
                                   ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => D1HSRXDATA(0),
      GlitchData                => D1HSRXDATA_GlitchData0,
      OutSignalName             => "D1HSRXDATA(0)",
      OutTemp                   => D1HSRXDATA_zd(0),
      Paths                     => ( 0 => (CKP_ipd'last_event,tpd_CKP_D1HSRXDATA_posedge(0) ,true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

	
      VitalPathDelay01 (
      OutSignal                 => D1HSRXDATA(1),
      GlitchData                => D1HSRXDATA_GlitchData1,
      OutSignalName             => "D1HSRXDATA(1)",
      OutTemp                   => D1HSRXDATA_zd(1),
      Paths                     => ( 0 => (CKP_ipd'last_event,tpd_CKP_D1HSRXDATA_posedge(1) ,true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => D1HSRXDATA(2),
      GlitchData                => D1HSRXDATA_GlitchData2,
      OutSignalName             => "D1HSRXDATA(2)",
      OutTemp                   => D1HSRXDATA_zd(2),
      Paths                     => ( 0 => (CKP_ipd'last_event,tpd_CKP_D1HSRXDATA_posedge(2) ,true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => D1HSRXDATA(3),
      GlitchData                => D1HSRXDATA_GlitchData3,
      OutSignalName             => "D1HSRXDATA(3)",
      OutTemp                   => D1HSRXDATA_zd(3),
      Paths                     => ( 0 => (CKP_ipd'last_event,tpd_CKP_D1HSRXDATA_posedge(3) ,true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => D1HSRXDATA(4),
      GlitchData                => D1HSRXDATA_GlitchData4,
      OutSignalName             => "D1HSRXDATA(4)",
      OutTemp                   => D1HSRXDATA_zd(4),
      Paths                     => ( 0 => (CKP_ipd'last_event,tpd_CKP_D1HSRXDATA_posedge(4) ,true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => D1HSRXDATA(5),
      GlitchData                => D1HSRXDATA_GlitchData5,
      OutSignalName             => "D1HSRXDATA(5)",
      OutTemp                   => D1HSRXDATA_zd(5),
      Paths                     => ( 0 => (CKP_ipd'last_event,tpd_CKP_D1HSRXDATA_posedge(5) ,true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => D1HSRXDATA(6),
      GlitchData                => D1HSRXDATA_GlitchData6,
      OutSignalName             => "D1HSRXDATA(6)",
      OutTemp                   => D1HSRXDATA_zd(6),
      Paths                     => ( 0 => (CKP_ipd'last_event,tpd_CKP_D1HSRXDATA_posedge(6) ,true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => D1HSRXDATA(7),
      GlitchData                => D1HSRXDATA_GlitchData7,
      OutSignalName             => "D1HSRXDATA(7)",
      OutTemp                   => D1HSRXDATA_zd(7),
      Paths                     => ( 0 => (CKP_ipd'last_event,tpd_CKP_D1HSRXDATA_posedge(7) ,true)  ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);


      VitalPathDelay01 (
      OutSignal                 => D1SYNC,
      GlitchData                => D1SYNC_GlitchData,
      OutSignalName             => "D1SYNC",
      OutTemp                   => D1SYNC_zd,
      Paths                     => ( 0 => (CKP_ipd'last_event, tpd_CKP_D1SYNC_posedge, true)),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);


      VitalPathDelay01 (
      OutSignal                 => D1ERRSYNC,
      GlitchData                => D1ERRSYNC_GlitchData,
      OutSignalName             => "D1ERRSYNC",
      OutTemp                   => D1ERRSYNC_zd,
      Paths                     => ( 0 => (CKP_ipd'last_event, tpd_CKP_D1ERRSYNC_posedge, true)),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

      VitalPathDelay01 (
      OutSignal                 => D1NOSYNC,
      GlitchData                => D1NOSYNC_GlitchData,
      OutSignalName             => "D1NOSYNC",
      OutTemp                   => D1NOSYNC_zd,
      Paths                     => ( 0 => (CKP_ipd'last_event, tpd_CKP_D1NOSYNC_negedge, true)),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);


      VitalPathDelay01 (
      OutSignal                 => CLKDRXLPP,
      GlitchData                => CLKDRXLPP_GlitchData,
      OutSignalName             => "CLKDRXLPP",
      OutTemp                   => CLKDRXLPP_zd,
      Paths                     => ( 0 => (CKP_ipd'last_event, tpd_CKP_CLKDRXLPP, true)
                                   ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);


      VitalPathDelay01 (
      OutSignal                 => CLKDRXLPN,
      GlitchData                => CLKDRXLPN_GlitchData,
      OutSignalName             => "CLKDRXLPN",
      OutTemp                   => CLKDRXLPN_zd,
      Paths                     => ( 0 => (CKN_ipd'last_event, tpd_CKN_CLKDRXLPN, true)
                                   ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);


      VitalPathDelay01 (
      OutSignal                 => CLKHSBYTE,
      GlitchData                => CLKHSBYTE_GlitchData,
      OutSignalName             => "CLKHSBYTE",
      OutTemp                   => CLKHSBYTE_zd,
      Paths                     => ( 0 => (CKP_ipd'last_event, tpd_CKP_CLKHSBYTE, true)
                                   ),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
end process VITALPathDelay;
	
end SB_MIPI_RX_2LANE_V; 


----------------------------------------------------------------------------------
-- 			SF16K DEVICE PRIMITIVES 				--		
-- 	# SB_MAC16	# SB_IO_DLY	# SB_MIPI_TX_4LANE	#16K BRAM   	--
----------------------------------------------------------------------------------

---------------------------------------------------------------------------
----			 	REG_BYPASS_MUX  			---	
---------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;

entity REG_BYPASS_MUX is 
  	generic ( 
		DATA_WIDTH : integer 		 := 16 ) ; 
	port 	(
		CLK	   : in std_logic ; 
		RST 	   : in std_logic; 
		ENA	   : in std_logic ;
		D	   : in  std_logic_vector(DATA_WIDTH-1 downto 0);
		SELM	   : in std_logic ;
		Q          : out  std_logic_vector(DATA_WIDTH-1	downto 0)  
		); 
end REG_BYPASS_MUX; 

architecture REG_BYPASS_MUX_ARCH of REG_BYPASS_MUX is 

  signal REG_INTERNAL : std_logic_vector(DATA_WIDTH-1 downto 0); 
	
begin 

 dffe_proc: process(CLK,RST,ENA) 
 begin 
	 if (RST = '1') then 
		REG_INTERNAL <= (others => '0'); 
	 elsif rising_edge(CLK) then 
		if (ENA ='1') then
			REG_INTERNAL <= D ;
   	 	else  
			REG_INTERNAL <= REG_INTERNAL ; 
		end if; 	
	end if; 
 end process dffe_proc; 

 
 dataselmux_proc: process(SELM,REG_INTERNAL,D) 
 begin 
 	case SELM is 
	when '0' => Q <= D; 
	when '1' =>  Q<=REG_INTERNAL; 
	when others =>  Q<=(others =>'0'); 
	end case; 
 end process dataselmux_proc; 		
		 
end  REG_BYPASS_MUX_ARCH; 


---------------------------------------------------------------------------
----			 	ha		  			---	
---------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;

entity ha is
	port (
		 A	: in 	std_logic ; 
		 B	: in	std_logic ; 
		 Sum	: out 	std_logic ; 
		 Cout   : out 	std_logic  
	       );

end ha; 


architecture ha_arch of ha is 
begin 
	Cout <= A and  B;
	Sum  <= A xor  B;

end ha_arch;

---------------------------------------------------------------------------
----			 	fa		  			---	
---------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;


entity fa is
	port (
		 A	: in 	std_logic ; 
		 B	: in	std_logic ;
		 C	: in 	std_logic ; 
		 Sum	: out 	std_logic ; 
		 Cout   : out 	std_logic  
	       );

end fa; 


architecture fa_arch of fa is 
begin 
	 Cout <= not ((not(A and B)) and  (not(B and C)) and (not(A and C)));
	 Sum  <= A xor B xor C;

end fa_arch; 

-----------------------------------------------------------------------------
------			 	mpfa 		  			---	
---------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;


entity mpfa  is 
	port ( 
		A 	: in 	std_logic ; 
		B	: in	std_logic ;	
		Cin	: in	std_logic ; 
	        Sum	: out 	std_logic ;
		p	: out	std_logic ; 			
		g_b	: out 	std_logic 
	     ); 

end mpfa; 

architecture mpfa_arch of mpfa  is 
   signal p_temp : std_logic;  	
begin 
	 p_temp   <= A xor B;
	
	 g_b <= not(A and B);
  	 p   <= p_temp; 	
	 Sum <= p_temp xor Cin;


end mpfa_arch ; 


-----------------------------------------------------------------------------
----			 	mclg4 		  			---	
---------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;

entity  mclg4 is 
	port ( 
	     	g_b 	: in 	std_logic_vector( 3 downto 0 ) ; 	
	 	p	: in 	std_logic_vector( 3 downto 0 ) ;
		cin	: in 	std_logic ; 
		g_o	: out	std_logic ; 
		p_o	: out 	std_logic ; 
		cout	: out	std_logic_vector ( 3 downto 0 ) 	
		); 
end mclg4; 

architecture mclg4_arch of mclg4 is 

 signal 	s1, s2, s3, s4, s5, s6,s7,s8,s9 : std_logic ;
 signal 	g : std_logic_vector( 2 downto 0 ) ;

begin 

	g(0) <= not(g_b(0));
	g(1) <= not(g_b(1));
	g(2) <= not(g_b(2));

	cout(0) <= '0';		-- Added to remove warning.  
	s1   <= not(p(0) and  cin);
	cout(1)  <= not (g_b(0) and  s1);

	s2 <= not (p(1) and g(0));
	s3 <= not (p(1) and  p(0) and  cin);
	cout(2) <= not(g_b(1) and s2 and  s3);

	s4 <= not(p(2) and  g(1));
	s5 <= not (p(2) and  p(1)  and  g(0));
	s6 <= not(p(2) and p(1) and  p(0) and  cin);
	cout(3) <= not (g_b(2) and  s4 and  s5 and s6);

	s7 <= not(p(3) and  g(2));
	s8 <= not(p(3) and  p(2) and  g(1));
	s9 <= not(p(3) and  p(2) and  p(1) and  g(0));
	g_o <= not(g_b(3) and  s7 and s8 and s9);

	p_o <=(p(3) and  p(2) and  p(1) and  p(0));

end mclg4_arch; 


---------------------------------------------------------------------------
----			 	mclg16 		  			---	
---------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;


entity  mclg16 is 
	port ( 
		g 	: in 	std_logic_vector( 3 downto 0) ; 
		p	: in	std_logic_vector( 3 downto 0) ; 
		cin	: in	std_logic ;
	  	g_o	: out	std_logic ; 
		p_o	: out	std_logic ; 
		cout	: out	std_logic_vector( 3 downto 0) 
 	     ); 
			
end mclg16;

architecture mclg16_arch of mclg16 is 

  signal s1, s2, s3, s4, s5, s6, s7,s8,s9 : std_logic ;

begin 


	cout(0) <= '0';		-- Added to remove warning.  

	s1 <= not( p(0) and  cin );
	cout(1) <= not( not(g(0)) and  s1 );

	s2 <= not ( p(1) and  g(0) );
	s3 <= not ( p(1) and  p(0) and  cin );
	cout(2) <= not ( not(g(1)) and  s2 and  s3 );

	s4 <= not( p(2) and  g(1) );
	s5 <= not( p(2) and p(1) and g(0) );
	s6 <= not( p(2) and p(1) and  p(0) and  cin );
	cout(3) <= not( not( g(2) ) and  s4 and  s5 and  s6 );

	s7 <= not ( p(3) and  g(2));
	s8 <= not ( p(3) and  p(2) and  g(1) );
	s9 <= not ( p(3) and  p(2) and  p(1) and  g(0) );
	g_o <= not( not(g(3)) and  s7 and  s8 and  s9 );

	p_o <= ( p(3) and  p(2) and p(1) and  p(0) );

end mclg16_arch; 

-------------------------------------------------------------------------
--			 fcla16			  			---	
---------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;

entity  fcla16 is 
	port  (	
		Sum	: out 	std_logic_vector( 15 downto 0); 
	        G	: out 	std_logic ; 
		P	: out 	std_logic ; 
		A	: in	std_logic_vector( 15 downto 0 );
		B	: in 	std_logic_vector( 15 downto 0 ); 
	 	Cin	: in 	std_logic
		);
end fcla16; 


architecture fcla16_arch of fcla16 is 

 component mpfa  is
        port (
                A       : in    std_logic ;
                B       : in    std_logic ;
                Cin     : in    std_logic ;
                Sum     : out   std_logic ;
                p       : out   std_logic ;
                g_b     : out   std_logic
             );
 end component;

 component mclg4 is
        port (
                g_b     : in    std_logic_vector( 3 downto 0 ) ;
                p       : in    std_logic_vector( 3 downto 0 ) ;
                cin     : in    std_logic ;
                g_o     : out   std_logic ;
                p_o     : out   std_logic ;
                cout    : out   std_logic_vector ( 3 downto 0 )
                );
 end component;
 
 component  mclg16 is 
	port ( 
		g 	: in 	std_logic_vector( 3 downto 0) ; 
		p	: in	std_logic_vector( 3 downto 0) ; 
		cin	: in	std_logic ;
	  	g_o	: out	std_logic ; 
		p_o	: out	std_logic ; 
		cout	: out	std_logic_vector( 3 downto 0) 
 	     ); 
 end component;
 
 signal  gtemp1_b : std_logic_vector( 15 downto 0);
 signal ptemp1 	: std_logic_vector (15 downto 0) ;
 signal ctemp1 	: std_logic_vector (15 downto 0) ;

 signal ctemp2  : std_logic_vector ( 3 downto 0) ;
 signal  gouta 	: std_logic_vector ( 3 downto 0) ; 
 signal  pouta 	: std_logic_vector ( 3 downto 0) ;

begin 

 r01 : mpfa port map (g_b => gtemp1_b(0), p=>ptemp1(0), Sum=>Sum(0), A=>A(0), B=>B(0), Cin=>Cin      );
 r02 : mpfa port map (g_b => gtemp1_b(1), p=>ptemp1(1), Sum=>Sum(1), A=>A(1), B=>B(1), Cin=>ctemp1(1) );
 r03 : mpfa port map (g_b =>gtemp1_b(2), p=>ptemp1(2), Sum=>Sum(2), A=>A(2), B=>B(2), Cin=>ctemp1(2)  );
 r04 : mpfa port map (g_b => gtemp1_b(3), p=>ptemp1(3), Sum=>Sum(3), A=>A(3), B=>B(3), Cin=>ctemp1(3) );
 b1  : mclg4 port map (cout=>ctemp1(3 downto 0), g_o=>gouta(0), p_o=>pouta(0), g_b=>gtemp1_b(3 downto 0),p=>ptemp1(3 downto 0), cin=>Cin );

 r05 : mpfa port map (g_b=>gtemp1_b(4), p=>ptemp1(4), Sum=>Sum(4), A=>A(4), B=>B(4), Cin=>ctemp2(1) );
 r06 : mpfa port map (g_b=>gtemp1_b(5), p=>ptemp1(5), Sum=>Sum(5), A=>A(5), B=>B(5), Cin=>ctemp1(5) );
 r07 : mpfa port map (g_b=>gtemp1_b(6), p=>ptemp1(6), Sum=>Sum(6), A=>A(6), B=>B(6), Cin=>ctemp1(6) );
 r08 : mpfa port map (g_b=>gtemp1_b(7), p=>ptemp1(7), Sum=>Sum(7), A=>A(7), B=>B(7), Cin=>ctemp1(7) );
 b2  : mclg4 port map (cout=>ctemp1(7 downto 4), g_o=>gouta(1), p_o=>pouta(1), g_b=>gtemp1_b(7 downto 4), p=>ptemp1(7 downto 4), cin=>ctemp2(1) );

 r09 : mpfa port map (g_b=>gtemp1_b(8), p=>ptemp1(8), Sum=>Sum(8), A=>A(8), B=>B(8), Cin=>ctemp2(2) );
 r10 : mpfa port map (g_b=>gtemp1_b(9), p=>ptemp1(9), Sum=>Sum(9), A=>A(9), B=>B(9), Cin=>ctemp1(9) );
 r11 : mpfa port map (g_b=>gtemp1_b(10), p=>ptemp1(10), Sum=>Sum(10), A=>A(10), B=>B(10), Cin=>ctemp1(10) );
 r12 : mpfa port map (g_b=>gtemp1_b(11), p=>ptemp1(11), Sum=>Sum(11), A=>A(11), B=>B(11), Cin=>ctemp1(11) );
 b3  : mclg4 port map (cout=>ctemp1(11 downto 8), g_o=>gouta(2), p_o=>pouta(2), g_b=>gtemp1_b(11 downto 8), p=>ptemp1(11 downto 8), cin=>ctemp2(2) );

 r13 : mpfa port map (g_b=>gtemp1_b(12), p=>ptemp1(12), Sum=>Sum(12), A=>A(12), B=>B(12), Cin=>ctemp2(3) );
 r14 : mpfa port map (g_b=>gtemp1_b(13), p=>ptemp1(13), Sum=>Sum(13), A=>A(13), B=>B(13), Cin=>ctemp1(13) );
 r15 : mpfa port map (g_b=>gtemp1_b(14), p=>ptemp1(14), Sum=>Sum(14), A=>A(14), B=>B(14), Cin=>ctemp1(14) );
 r16 : mpfa port map (g_b=>gtemp1_b(15), p=>ptemp1(15), Sum=>Sum(15), A=>A(15), B=>B(15), Cin=>ctemp1(15) );
 b4  : mclg4 port map (cout=>ctemp1(15 downto 12), g_o=>gouta(3), p_o=>pouta(3), g_b=>gtemp1_b(15 downto 12), p=>ptemp1(15 downto 12), cin=>ctemp2(3) );

 b5  : mclg16 port map (cout=>ctemp2, g_o=>G, p_o=>P, g=>gouta, p=>pouta, cin=>Cin );

end fcla16_arch; 


---------------------------------------------------------------------------
--			  fcla8	 		  			---	
---------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;


entity fcla8 is 
	port 
	  (
		Sum 	: out 	std_logic_vector( 7 downto 0); 
		G	: out 	std_logic ; 
		P	: out 	std_logic ;
		A	: in	std_logic_vector( 7 downto 0);  
		B	: in 	std_logic_vector( 7 downto 0); 
		Cin     : in	std_logic 
	  );
end fcla8; 

architecture fcla8_arch of fcla8 is 

  component mpfa  is
        port (
                A       : in    std_logic ;
                B       : in    std_logic ;
                Cin     : in    std_logic ;
                Sum     : out   std_logic ;
                p       : out   std_logic ;
                g_b     : out   std_logic
             );
 end component;

 component mclg4 is
        port (
                g_b     : in    std_logic_vector( 3 downto 0 ) ;
                p       : in    std_logic_vector( 3 downto 0 ) ;
                cin     : in    std_logic ;
                g_o     : out   std_logic ;
                p_o     : out   std_logic ;
                cout    : out   std_logic_vector ( 3 downto 0 )
                );
 end component ;


 signal	gtemp1	: std_logic_vector( 7 downto 0) ;
 signal	ptemp1	: std_logic_vector( 7 downto 0) ;
 signal	ctemp1	: std_logic_vector( 7 downto 0) ;
 signal	ctemp2	: std_logic ; 
 signal	gouta	: std_logic_vector( 1 downto 0) ;
 signal	pouta	: std_logic_vector( 1 downto 0) ;

begin 


 r01 : mpfa port map  (g_b=>gtemp1(0), p=>ptemp1(0), Sum=>Sum(0), A=>A(0), B=>B(0), Cin=>Cin );
 r02 : mpfa port map (g_b=>gtemp1(1), p=>ptemp1(1), Sum=>Sum(1), A=>A(1), B=>B(1), Cin=>ctemp1(1) );
 r03 : mpfa port map (g_b=>gtemp1(2), p=>ptemp1(2), Sum=>Sum(2), A=>A(2), B=>B(2), Cin=>ctemp1(2) );
 r04 : mpfa port map (g_b=>gtemp1(3), p=>ptemp1(3), Sum=>Sum(3), A=>A(3), B=>B(3), Cin=>ctemp1(3) );
 b1  : mclg4 port map (cout=>ctemp1(3 downto 0), g_o=>gouta(0), p_o=>pouta(0), g_b=>gtemp1( 3 downto 0), p=>ptemp1(3 downto 0), cin=>Cin );

 r05 : mpfa port map (g_b=>gtemp1(4), p=>ptemp1(4), Sum=>Sum(4), A=>A(4), B=>B(4), Cin=>ctemp2 );
 r06 : mpfa port map (g_b=>gtemp1(5), p=>ptemp1(5), Sum=>Sum(5), A=>A(5), B=>B(5), Cin=>ctemp1(5) );
 r07 : mpfa port map (g_b=>gtemp1(6), p=>ptemp1(6), Sum=>Sum(6), A=>A(6), B=>B(6), Cin=>ctemp1(6) );
 r08 : mpfa port map (g_b=>gtemp1(7), p=>ptemp1(7), Sum=>Sum(7), A=>A(7), B=>B(7), Cin=>ctemp1(7));
 b2  : mclg4 port map (cout=>ctemp1(7 downto 4), g_o=>gouta(1), p_o=>pouta(1), g_b=>gtemp1(7 downto 4), p=>ptemp1(7 downto 4), cin=>ctemp2 );

 ctemp2 <= not( not(gouta(0)) and not(pouta(0) and  Cin ));

 G <= not( ( not (gouta(1)) ) and ( not (pouta(1) and  gouta(0)) ) );
 P <= pouta(1) and  pouta(0);

end fcla8_arch ; 


---------------------------------------------------------------------------
----			ADDER_A_IN_MUX 		  			---	
---------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;

entity ADDER_A_IN_MUX is 
	port  (
		ACCUMULATOR_REG  	: in std_logic_vector(15 downto 0); 
		DIRECT_INPUT		: in std_logic_vector(15 downto 0); 
		SELM 			: in std_logic ;
		ADDER_A_MUX		: out std_logic_vector( 15 downto 0) 
	        );
end ADDER_A_IN_MUX ; 


architecture ADDER_A_IN_MUX_ARCH of ADDER_A_IN_MUX is 
begin

	process(SELM , DIRECT_INPUT , ACCUMULATOR_REG) is 
	begin 
		case (SELM) is 
		when '0'    => ADDER_A_MUX <= ACCUMULATOR_REG;  
		when '1'    => ADDER_A_MUX <= DIRECT_INPUT; 
		when others => ADDER_A_MUX <= (others => 'X'); 
		end case;
	end process; 

end ADDER_A_IN_MUX_ARCH; 


---------------------------------------------------------------------------
----			  ADDER_B_IN_MUX	  			---	
---------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;


entity  ADDER_B_IN_MUX  is 
	port (
		MULT_INPUT  	: in 	std_logic_vector( 15 downto 0 ); 
		MULT_8x8 	: in 	std_logic_vector( 15 downto 0 ); 
		MULT_16x16 	: in	std_logic_vector( 15 downto 0 ); 
		SIGNEXTIN 	: in	std_logic ; 
		SELM 		: in 	std_logic_vector ( 1 downto 0) ;
		ADDER_B_MUX     : out   std_logic_vector ( 15 downto 0)
	       );
end ADDER_B_IN_MUX ; 



architecture ADDER_B_IN_MUX_ARCH of ADDER_B_IN_MUX is 
begin 
	
 process (SELM , MULT_INPUT , MULT_8x8 , MULT_16x16 , SIGNEXTIN) is 
 begin 	
      case(SELM) is
        when "00" => ADDER_B_MUX <= MULT_INPUT ; 
        when "01" => ADDER_B_MUX <= MULT_8x8 ; 
        when "10" => ADDER_B_MUX <= MULT_16x16; 
	when "11" => ADDER_B_MUX <=(others => SIGNEXTIN );
	when others => ADDER_B_MUX <= (others => 'X');  
      end case ;
  end process; 	
	
end ADDER_B_IN_MUX_ARCH;  


-----------------------------------------------------------------------------
----			  CARRY_IN_MUX		  			---	
---------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;

entity  CARRY_IN_MUX is 
	port (
		CICAS		: in std_logic ; 
		CI		: in std_logic ; 
		CARRYMUX_SEL 	: in std_logic_vector( 1 downto 0); 
		ADDER_CI	: out std_logic 
	   );
end CARRY_IN_MUX;

architecture CARRY_IN_MUX_ARCH of CARRY_IN_MUX is  	
begin 
	
 process(CARRYMUX_SEL, CICAS ,CI) is 
 begin 	
      case(CARRYMUX_SEL) is 
         when "00" =>  ADDER_CI <= '0' ; 
         when "01" =>  ADDER_CI <= '1' ; 
         when "10" =>  ADDER_CI <= CICAS; 
         when "11" =>  ADDER_CI <= CI; 
	when others => ADDER_CI <= '0'; 
      end case; 	 
  end process;

end CARRY_IN_MUX_ARCH; 

	
-------------------------------------------------------------------------------
-----			OUT_MUX_4   		  			---	
---------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;

entity OUT_MUX_4 is 
	port (
		ADDER_COMBINATORIAL  	: in std_logic_vector( 15 downto 0); 
	    	ACCUM_REGISTER 		: in std_logic_vector( 15 downto 0);
		MULT_8x8 		: in std_logic_vector( 15 downto 0); 
		MULT_16x16 		: in std_logic_vector( 15 downto 0);
		SELM 			: in std_logic_vector( 1 downto 0);
		OUT_O  			: out std_logic_vector( 15 downto 0)	
	 ) ;

end  OUT_MUX_4; 

architecture OUT_MUX_4_ARCH of OUT_MUX_4 is 
begin 
	process (SELM, ADDER_COMBINATORIAL ,ACCUM_REGISTER , MULT_8x8 , MULT_16x16) is 
	begin 
		case (SELM) is 
         	when "00" => OUT_O <= ADDER_COMBINATORIAL ; 	-- Combinatorial Adder output.
         	when "01" => OUT_O <= ACCUM_REGISTER ; 		-- Accumulator register output.
	        when "10" => OUT_O <= MULT_8x8;  		--  MULT_8x8 output.  
         	when "11" => OUT_O <= MULT_16x16;  		--  MULT_16x16 output. 
	 	when others => OUT_O <= (others => 'X'); 	
      	end case;	 
	end process; 	

end OUT_MUX_4_ARCH; 


---------------------------------------------------------------------------
------			ACCUM_REG	  				---	
---------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;

entity  ACCUM_REG  is 
	port (
		D 	: in 	std_logic_vector ( 15 downto 0 ); 
		Q 	: out 	std_logic_vector ( 15 downto 0 ); 
		ENA 	: in	std_logic ; 
		CLK 	: in	std_logic ;
		RST     : in	std_logic 
	);

end ACCUM_REG; 


architecture ACCUM_REG_ARCH of ACCUM_REG is 
   
 signal Q_INTERNAL :  std_logic_vector ( 15 downto 0 ); 
 
begin 	
	process (CLK,RST,ENA) is 
	begin 
      		if (RST='1' ) then 		--  Syncronous reset overrides all other controls
			Q_INTERNAL <= (others => '0');
		elsif rising_edge (CLK) then 
		 	if (ENA ='1') then 			--  Update Q whenever LOAD or ENAble asserted
				Q_INTERNAL <=  D ;
			else
				Q_INTERNAL <= Q_INTERNAL ;
			end if; 
		end if; 
	end process ; 
	
	Q <= Q_INTERNAL; ---  after 1ns; 
	
end ACCUM_REG_ARCH;   


-----------------------------------------------------------------------------
----			LOAD_ADD_MUX   		  			---	
---------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;

entity LOAD_ADD_MUX is 
	port (
		ADDER_DATA	: in	std_logic_vector(15 downto 0); 	
		LOAD_DATA	: in   	std_logic_vector(15 downto 0); 
		LOAD		: in  	std_logic ; 	
		LDATAOUT	: out   std_logic_vector(15 downto 0)
  	      );
end LOAD_ADD_MUX; 

architecture LOAD_ADD_MUX_ARCH of LOAD_ADD_MUX is 
begin 
	process(LOAD, LOAD_DATA, ADDER_DATA) is 
	begin 
		case (LOAD) is 
		when '0' => LDATAOUT <= ADDER_DATA ; 
		when '1' => LDATAOUT <=LOAD_DATA ; 	
		when others => LDATAOUT <=(others => 'X'); 
		end case ; 	
	end process;  
	
end LOAD_ADD_MUX_ARCH; 

---------------------------------------------------------------------------
----			  ACCUM_ADDER 		  			---	
---------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;

entity  ACCUM_ADDER is 
	port  (
		A 	: in  	std_logic_vector ( 15  downto 0 ); 
		B 	: in 	std_logic_vector ( 15 downto 0 ); 
		ADDSUB 	: in	std_logic; 
		CI 	: in	std_logic ; 
		SUM 	: out 	std_logic_vector ( 15 downto 0 ); 
		COCAS 	: out 	std_logic ; 
		CO	: out   std_logic 
	       );

end ACCUM_ADDER; 

architecture ACCUM_ADDER_ARCH of ACCUM_ADDER is 

 component   fcla16 is
        port  (
                Sum     : out   std_logic_vector( 15 downto 0);
                G       : out   std_logic ;
                P       : out   std_logic ;
                A       : in    std_logic_vector( 15 downto 0 );
                B       : in    std_logic_vector( 15 downto 0 );
                Cin     : in    std_logic
                );
 end component;

 signal 	CLA16_g, CLA16_p : std_logic ;
 signal CLA16_SUM  : std_logic_vector ( 15 downto 0); 
 signal CLA16_A	  : std_logic_vector ( 15 downto 0);
 signal COCAS_temp : std_logic; 
 signal  j : integer;

begin 

 process(ADDSUB,COCAS_temp, A,CLA16_SUM) is 
 begin
	if (ADDSUB = '1') then 
		 CO <= not(COCAS_temp);
           for j in 0 to 15 loop  
		 CLA16_A(j) <= not( A(j));
		 SUM(j) <= not( CLA16_SUM(j));
	    end loop;
	else 
	   CO 			<= COCAS_temp;
	   CLA16_A(15 downto 0) <= A(15 downto 0);
	   SUM(15 downto 0) 	<= CLA16_SUM(15 downto 0);
	end if; 
 end process; 

 CLA16_ADDER  : fcla16 port map (
		Sum=>CLA16_SUM(15 downto 0),
		A=>CLA16_A(15 downto 0),
		B=>B(15 downto 0), 
		G=>CLA16_g,
		P=>CLA16_p,
		Cin=>CI );


  COCAS_temp <= not ( (not(CLA16_g)) and  (not(CLA16_p and CI)));
  COCAS      <= COCAS_temp; 	

end  ACCUM_ADDER_ARCH; 


---------------------------------------------------------------------------
----			MULT_ACCUM 		  			---	
---------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;

entity  MULT_ACCUM is 
	port  (
		DIRECT_INPUT	: in std_logic_vector ( 15 downto 0); 
		MULT_INPUT	: in std_logic_vector ( 15 downto 0);
    		MULT_8x8	: in std_logic_vector ( 15 downto 0);	
		MULT_16x16	: in std_logic_vector ( 15 downto 0);
		ADDSUB		: in std_logic ; 
		CLK		: in std_logic ;
    		CICAS		: in std_logic ;
    		CI		: in std_logic ;
		SIGNEXTIN	: in std_logic ;
		SIGNEXTOUT	: out std_logic ;
    		LDA		: in std_logic ; 
    		RST		: in std_logic ;
    		ENA		: in std_logic ;
    		COCAS		: out std_logic ;
    		CO		: out std_logic ;
    		O		: out std_logic_vector ( 15 downto 0);
		OUTMUX_SEL	: in std_logic_vector ( 1 downto 0);
		CARRYMUX_SEL	: in std_logic_vector ( 1 downto 0);
		ADDER_A_IN_SEL  : in std_logic;
		ADDER_B_IN_SEL  : in std_logic_vector ( 1 downto 0)
    		);

end MULT_ACCUM;

architecture MULT_ACCUM_ARCH of MULT_ACCUM is 

 component ADDER_A_IN_MUX is
        port  (
                ACCUMULATOR_REG         : in std_logic_vector(15 downto 0);
                DIRECT_INPUT            : in std_logic_vector(15 downto 0);
                SELM                    : in std_logic ;
                ADDER_A_MUX             : out std_logic_vector( 15 downto 0)
                );
 end component; 

 component  ADDER_B_IN_MUX  is
        port (
                MULT_INPUT      : in    std_logic_vector( 15 downto 0 );
                MULT_8x8        : in    std_logic_vector( 15 downto 0 );
                MULT_16x16      : in    std_logic_vector( 15 downto 0 );
                SIGNEXTIN       : in    std_logic ;
                SELM            : in    std_logic_vector ( 1 downto 0) ;
                ADDER_B_MUX     : out   std_logic_vector ( 15 downto 0)
               );
 end component; 

 component  CARRY_IN_MUX is
        port (
                CICAS           : in std_logic ;
                CI              : in std_logic ;
                CARRYMUX_SEL    : in std_logic_vector( 1 downto 0);
                ADDER_CI        : out std_logic
           );
 end component; 

 component OUT_MUX_4 is
        port (
                ADDER_COMBINATORIAL     : in std_logic_vector( 15 downto 0);
                ACCUM_REGISTER          : in std_logic_vector( 15 downto 0);
                MULT_8x8                : in std_logic_vector( 15 downto 0);
                MULT_16x16              : in std_logic_vector( 15 downto 0);
                SELM                    : in std_logic_vector( 1 downto 0);
                OUT_O                   : out std_logic_vector( 15 downto 0)
         ) ;

 end component;

 component  ACCUM_REG  is
        port (
                D       : in    std_logic_vector ( 15 downto 0 );
                Q       : out   std_logic_vector ( 15 downto 0 );
                ENA     : in    std_logic ;
                CLK     : in    std_logic ;
                RST     : in    std_logic
        );

 end component; 

 component LOAD_ADD_MUX is
        port (
                ADDER_DATA      : in    std_logic_vector(15 downto 0);
                LOAD_DATA       : in    std_logic_vector(15 downto 0);
                LOAD            : in    std_logic ;
                LDATAOUT        : out   std_logic_vector(15 downto 0)
              );
 end component; 

 component  ACCUM_ADDER is
        port  (
                A       : in    std_logic_vector ( 15  downto 0 );
                B       : in    std_logic_vector ( 15 downto 0 );
                ADDSUB  : in    std_logic;
                CI      : in    std_logic ;
                SUM     : out   std_logic_vector ( 15 downto 0 );
                COCAS   : out   std_logic ;
                CO      : out   std_logic
               );
 end component; 

  signal  ADDER_LOAD_MUX	: std_logic_vector ( 15 downto 0) ;
  signal  ACCUMULATOR_REG	: std_logic_vector ( 15 downto 0) ;
  signal  ADDER_SUM 		: std_logic_vector ( 15 downto 0) ;
  signal  ADDER_A_INPUT_MUX 	: std_logic_vector ( 15 downto 0) ;
  signal  ADDER_B_INPUT_MUX 	: std_logic_vector ( 15 downto 0) ;
  signal  ADDER_CI		: std_logic ; 

begin 
	 
 SIGNEXTOUT <= ADDER_B_INPUT_MUX(15);
  
 OUTPUT_MULTIPLEXER_TOP : OUT_MUX_4 port map (
		ADDER_COMBINATORIAL	=> ADDER_LOAD_MUX ,	
		ACCUM_REGISTER 		=> ACCUMULATOR_REG  ,
		MULT_8x8		=> MULT_8x8 ,
		MULT_16x16		=> MULT_16x16,
		SELM			=> OUTMUX_SEL(1 downto 0),
		OUT_O			=> O  
		 ) ;
 
 ACCUM_REG_TOP :  ACCUM_REG port map   (
		D	=> ADDER_LOAD_MUX,
		Q	=> ACCUMULATOR_REG ,
		ENA	=> ENA,
		CLK	=> CLK ,
		RST	=> RST
		);
	
 ACCUM_ADDER_TOP : ACCUM_ADDER port map (
		A	=> ADDER_A_INPUT_MUX,
		B	=> ADDER_B_INPUT_MUX,
		ADDSUB	=> ADDSUB,
		CI	=> ADDER_CI ,
		SUM	=> ADDER_SUM ,
		COCAS	=> COCAS,
		CO	=> CO
		);	

 LOAD_ADD_TOP : LOAD_ADD_MUX port map (
		ADDER_DATA	=> ADDER_SUM ,
		LOAD_DATA	=> DIRECT_INPUT,
		LOAD		=> LDA,
		LDATAOUT	=> ADDER_LOAD_MUX
		 );
 
 ADDER_A_IN_MUX_TOP : ADDER_A_IN_MUX port map  (
		ACCUMULATOR_REG	=> ACCUMULATOR_REG,
		DIRECT_INPUT	=> DIRECT_INPUT,
		SELM		=> ADDER_A_IN_SEL,
		ADDER_A_MUX	=> ADDER_A_INPUT_MUX
  		 );

 ADDER_B_IN_MUX_TOP : ADDER_B_IN_MUX port map (
   		MULT_INPUT	=> MULT_INPUT,
		MULT_8x8	=> MULT_8x8,
		MULT_16x16	=> MULT_16x16,
		SIGNEXTIN	=> SIGNEXTIN,
		SELM		=> ADDER_B_IN_SEL(1 downto 0),
		ADDER_B_MUX	=> ADDER_B_INPUT_MUX
		);	

 CARRY_IN_MUX_TOP : CARRY_IN_MUX port map (
		CICAS		=> CICAS ,
		CI		=> CI,
		CARRYMUX_SEL	=> CARRYMUX_SEL(1 downto 0),
		ADDER_CI	=> ADDER_CI
		);
	
end MULT_ACCUM_ARCH;  

---------------------------------------------------------------------------
----			booth_encoder		  			---	
---------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;


entity booth_encoder  is 
	port (	
		booth_single	:  out std_logic_vector(4 downto 0) ; 
		booth_double	:  out std_logic_vector(4 downto 0) ; 
		booth_negtive	:  out std_logic_vector(4 downto 0) ; 
		multiplier	:  in std_logic_vector(7 downto 0) ; 
		signed_mpy	:  in std_logic 
	    );
end booth_encoder; 

architecture booth_encoder_arch of booth_encoder is 
 signal booth_in 	:  std_logic_vector(10 downto 0);
 signal sign_ext   :  std_logic_vector( 1 downto 0);
begin 

	process(signed_mpy, multiplier) is  
	begin 
	case(signed_mpy) is 
	when '0' =>  sign_ext <= "00"; 
	when '1'  => sign_ext <= multiplier(7) & multiplier(7) ;  
	when others => sign_ext <=(others => '0'); 
	end case; 
	end process; 	
	
	  booth_in <= sign_ext & multiplier(7 downto 0) & '0';

	  booth_negtive(0) <= booth_in(2);
	  booth_negtive(1) <= booth_in(4);
	  booth_negtive(2) <= booth_in(6);
	  booth_negtive(3) <= booth_in(8);
	  booth_negtive(4) <= booth_in(10);

	  booth_single(0) <= booth_in(0) xor booth_in(1);
	  booth_single(1) <= booth_in(2) xor booth_in(3);
	  booth_single(2) <= booth_in(4) xor booth_in(5);
	  booth_single(3) <= booth_in(6) xor booth_in(7);
	  booth_single(4) <= booth_in(8) xor booth_in(9);

	  booth_double(0)<= not( not( booth_in(0) and booth_in(1) and  not( booth_in(2)) ) and  not( not( booth_in(0)) and  not( booth_in(1)) and booth_in(2)));
	  booth_double(1)<= not( not( booth_in(2) and booth_in(3) and  not( booth_in(4)) ) and  not( not( booth_in(2)) and  not( booth_in(3)) and booth_in(4)));
	  booth_double(2)<= not( not( booth_in(4) and booth_in(5) and  not( booth_in(6)) ) and  not( not( booth_in(4)) and  not( booth_in(5)) and booth_in(6)));
	  booth_double(3)<= not( not( booth_in(6) and booth_in(7) and  not( booth_in(8)) ) and  not( not( booth_in(6)) and  not( booth_in(7)) and booth_in(8)));
	  booth_double(4)<= not( not( booth_in(8) and booth_in(9) and  not( booth_in(10))) and  not( not( booth_in(8)) and  not( booth_in(9)) and booth_in(10)));

end booth_encoder_arch; 



---------------------------------------------------------------------------
----			booth_selector 		  			---	
---------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;

entity  booth_selector is 
	port 	(
		pp_out		: out std_logic_vector(44 downto 0); 
		booth_single 	: in  std_logic_vector(4 downto 0); 
		booth_double    : in std_logic_vector(4 downto 0);
		booth_negtive   : in std_logic_vector(4 downto 0); 
		multiplicand    : in std_logic_vector(7 downto 0);
		signed_mpy      : in std_logic 
		);
end booth_selector; 


architecture booth_selector_arch of booth_selector is 

 signal j 		    : integer ;
 signal pp0,pp1,pp2,pp3,pp4 : std_logic_vector ( 8 downto 0);
 signal bs_in 		    : std_logic_vector ( 9 downto 0);
 signal sign_ext	    : std_logic;

begin 

	process(signed_mpy,multiplicand) is
        begin
        case(signed_mpy) is
	        when '0' =>  sign_ext <= '0';
        	when '1'  => sign_ext <= multiplicand(7) ; 
	       when others => sign_ext <= '0';
        end case;
        end process;

	pp_out <= pp4 & pp3 & pp2 & pp1 &  pp0; 


	bs_in <=sign_ext & multiplicand(7 downto 0) & '0';

	process (booth_negtive, booth_single , bs_in , booth_double)
	begin
	for j in 0 to 8  loop 
		pp0(j) <= (booth_negtive(0) xor not(not(booth_single(0) and bs_in(j+1)) and  not(booth_double(0) and  bs_in(j))) );
		pp1(j) <= (booth_negtive(1) xor not(not(booth_single(1) and  bs_in(j+1)) and  not(booth_double(1) and  bs_in(j))));
		pp2(j) <= (booth_negtive(2) xor not(not(booth_single(2) and bs_in(j+1)) and not(booth_double(2) and bs_in(j))));
		pp3(j) <= (booth_negtive(3) xor not(not(booth_single(3) and bs_in(j+1)) and not(booth_double(3) and bs_in(j))));
		pp4(j) <= (booth_negtive(4) xor not(not(booth_single(4) and bs_in(j+1)) and not(booth_double(4) and bs_in(j))));
	end loop; 
	end process;  

end  booth_selector_arch; 


---------------------------------------------------------------------------
----			MPY8x8 	 	  			---	
---------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;

entity MPY8x8 is 
	port 	(
		csa_a		: out std_logic_vector( 15 downto 0); 
		csa_b		: out std_logic_vector( 15 downto 0);
		multiplicand    : in  std_logic_vector( 7 downto 0);
		multiplier      : in  std_logic_vector( 7 downto 0); 
		signed_MPD      : std_logic ;    
		signed_MPR      : std_logic
		);
end MPY8x8; 

architecture MPY8x8_ARCH of MPY8x8 is 

 component booth_encoder  is
        port (
                booth_single    :  out std_logic_vector(4 downto 0) ;
                booth_double    :  out std_logic_vector(4 downto 0) ;
                booth_negtive   :  out std_logic_vector(4 downto 0) ;
                multiplier      :  in std_logic_vector(7 downto 0) ;
                signed_mpy      :  in std_logic
            );
 end component;

 component booth_selector is 
	port 	(
		pp_out		: out std_logic_vector(44 downto 0); 
		booth_single 	: in  std_logic_vector(4 downto 0); 
		booth_double    : in std_logic_vector(4 downto 0);
		booth_negtive   : in std_logic_vector(4 downto 0); 
		multiplicand    : in std_logic_vector(7 downto 0);
		signed_mpy      : in std_logic 
		);
 end component;

 component ha is
        port (
                 A      : in    std_logic ;
                 B      : in    std_logic ;
                 Sum    : out   std_logic ;
                 Cout   : out   std_logic
               );

 end component;

 component fa is
        port (
                 A      : in    std_logic ;
                 B      : in    std_logic ;
                 C      : in    std_logic ;
                 Sum    : out   std_logic ;
                 Cout   : out   std_logic
               );

 end component;

 signal	booth_single		: std_logic_vector( 4 downto 0) ;
 signal	booth_double       	: std_logic_vector( 4 downto 0) ; 
 signal	booth_negtive      	: std_logic_vector( 4 downto 0) ;
 signal	pp_sign            	: std_logic_vector( 4 downto 0) ;
 signal	pp_out            	: std_logic_vector( 44 downto 0) ;
 signal	PP0,PP1,PP2,PP3,PP4 	: std_logic_vector( 8 downto 0) ; 
 
 signal current_MPD_sign	: std_logic ; 


 signal j : integer ; 
 signal  booth_single_b, booth_double_b, booth_negtive_b :  std_logic_vector( 4 downto 0);

  --- WCSA step#1 Signals  
  signal	FA1_R00C14_C, FA1_R00C14_S: std_logic;
  signal	FA1_R00C13_C, FA1_R00C13_S: std_logic;
  signal	FA1_R00C12_C, FA1_R00C12_S: std_logic;
  signal	FA1_R00C11_C, FA1_R00C11_S: std_logic;
  signal	HA1_R03C11_C, HA1_R03C11_S: std_logic;
  signal	FA1_R00C10_C, FA1_R00C10_S: std_logic;
  signal	HA1_R03C10_C, HA1_R03C10_S: std_logic;
  signal	FA1_R00C09_C, FA1_R00C09_S: std_logic;
  signal	HA1_R03C09_C, HA1_R03C09_S: std_logic;
  signal	FA1_R00C08_C, FA1_R00C08_S: std_logic;
  signal	FA1_R03C08_C, FA1_R03C08_S: std_logic;
  signal	FA1_R00C07_C, FA1_R00C07_S: std_logic;
  signal	FA1_R00C06_C, FA1_R00C06_S: std_logic;
  signal	HA1_R03C06_C, HA1_R03C06_S: std_logic;
  signal	FA1_R00C05_C, FA1_R00C05_S: std_logic;
  signal	FA1_R00C04_C, FA1_R00C04_S: std_logic;
  signal	FA1_R00C02_C, FA1_R00C02_S: std_logic;
  
  --- WCSA step#2 Signals 
  signal	FA2_R00C15_C, FA2_R00C15_S: std_logic;
  signal	HA2_R00C14_C, HA2_R00C14_S: std_logic;
  signal	HA2_R00C13_C, HA2_R00C13_S: std_logic;
  
  signal	FA2_R00C12_C, FA2_R00C12_S: std_logic;
  signal	FA2_R00C11_C, FA2_R00C11_S: std_logic;
  signal	FA2_R00C10_C, FA2_R00C10_S: std_logic;
  signal	FA2_R00C09_C, FA2_R00C09_S: std_logic;
  signal	FA2_R00C08_C, FA2_R00C08_S: std_logic;
  signal	FA2_R00C07_C, FA2_R00C07_S: std_logic;
  signal	FA2_R00C06_C, FA2_R00C06_S: std_logic;
  
  signal	FA2_R00C03_C, FA2_R00C03_S: std_logic;
  
  -- WCSA step#3 Signals 
  signal	HA3_R00C15_C, HA3_R00C15_S: std_logic;
  signal	HA3_R00C14_C, HA3_R00C14_S: std_logic;
  signal	HA3_R00C13_C, HA3_R00C13_S: std_logic;
  signal	FA3_R00C12_C, FA3_R00C12_S: std_logic;
  signal	FA3_R00C11_C, FA3_R00C11_S: std_logic;
  signal	FA3_R00C10_C, FA3_R00C10_S: std_logic;
  signal	FA3_R00C09_C, FA3_R00C09_S: std_logic;
  
  signal	HA3_R00C08_C, HA3_R00C08_S: std_logic;
  signal	FA3_R00C07_C, FA3_R00C07_S: std_logic;
  
  signal	HA3_R00C05_C, HA3_R00C05_S: std_logic;
  signal	FA3_R00C04_C, FA3_R00C04_S: std_logic;
 

 signal 	pp_sign_2_not, pp_sign_0_not 	: std_logic ; 
 signal 	pp_sign_1_not, pp_sign_3_not	: std_logic ; 
 

begin
 
 PP0 <= pp_out(8 downto 0); 
 PP1 <= pp_out(17 downto 9); 
 PP2 <= pp_out(26 downto 18); 
 PP3 <= pp_out(35 downto 27); 
 PP4 <= pp_out(44 downto 36); 
 --
 booth_encoder_i :  booth_encoder port map (
		booth_single	=>booth_single, 
		booth_double	=>booth_double, 
		booth_negtive	=>booth_negtive, 
		multiplier	=>multiplier,
		signed_mpy	=>signed_MPR
		);

 booth_selector_i :  booth_selector port map (
		pp_out 		=> pp_out,
		booth_single	=> booth_single, 
		booth_double 	=> booth_double, 
		booth_negtive	=> booth_negtive,
		multiplicand	=> multiplicand,
		signed_mpy	=>signed_MPD
		);

 current_MPD_sign <= multiplicand(7) and  signed_MPD;

 process(booth_single, booth_double,booth_negtive)
 begin
 	for j in 0 to 4 loop 
		    booth_single_b(j) <=not(booth_single(j));
	            booth_double_b(j) <=not(booth_double(j));
	            booth_negtive_b(j) <= not(booth_negtive(j));
	end loop ; 			
 end process; 

  --
	 pp_sign(0) <= ((booth_negtive(0) xor  current_MPD_sign) and (not(booth_single_b(0) and  booth_double_b(0) and  booth_negtive_b(0)))) or ( booth_single_b(0) and  booth_double_b(0) and  booth_negtive(0) ) ;
	 pp_sign(1) <= ((booth_negtive(1) xor  current_MPD_sign) and (not(booth_single_b(1) and  booth_double_b(1) and  booth_negtive_b(1)))) or (booth_single_b(1) and  booth_double_b(1) and  booth_negtive(1));
	 pp_sign(2) <= ((booth_negtive(2) xor  current_MPD_sign) and (not(booth_single_b(2) and  booth_double_b(2) and  booth_negtive_b(2)))) or (booth_single_b(2) and  booth_double_b(2) and  booth_negtive(2));
	 pp_sign(3) <= ((booth_negtive(3) xor  current_MPD_sign) and (not(booth_single_b(3) and  booth_double_b(3) and  booth_negtive_b(3)))) or (booth_single_b(3) and  booth_double_b(3) and  booth_negtive(3));
	 pp_sign(4) <= ((booth_negtive(4) xor  current_MPD_sign) and (not(booth_single_b(4) and  booth_double_b(4) and  booth_negtive_b(4)))) or (booth_single_b(4) and  booth_double_b(4) and booth_negtive(4));

  -- WCSA step#1

  pp_sign_0_not <= not(pp_sign(0));  
  pp_sign_1_not <= not(pp_sign(1));	
  pp_sign_2_not <= not(pp_sign(2));
  pp_sign_3_not <= not(pp_sign(3));
  	
  FA1_R00C14 : fa port map (Cout=>FA1_R00C14_C, Sum=>FA1_R00C14_S, A=>'1', B=>PP3(8), C=>PP4(6) );
  FA1_R00C13 : fa port map (Cout=>FA1_R00C13_C, Sum=>FA1_R00C13_S, A=>pp_sign_2_not , B=>PP3(7), C=>PP4(5) );
  FA1_R00C12 : fa port map (Cout=>FA1_R00C12_C, Sum=>FA1_R00C12_S, A=>'1', B=>PP2(8), C=>PP3(6) );
  FA1_R00C11 : fa port map (Cout=>FA1_R00C11_C, Sum=>FA1_R00C11_S, A=>pp_sign_0_not , B=>pp_sign_1_not, C=>PP2(7) );
  HA1_R03C11 : ha port map (Cout=>HA1_R03C11_C, Sum=>HA1_R03C11_S, A=>PP3(5), B=>PP4(3) );

  FA1_R00C10 : fa port map (Cout=>FA1_R00C10_C, Sum=>FA1_R00C10_S, A=>pp_sign(0), B=>PP1(8), C=>PP2(6) );
  HA1_R03C10 : ha port map (Cout=>HA1_R03C10_C, Sum=>HA1_R03C10_S, A=>PP3(4), B=>PP4(2) );

  FA1_R00C09 : fa port map (Cout=>FA1_R00C09_C, Sum=>FA1_R00C09_S, A=>pp_sign(0), B=>PP1(7) , C=>PP2(5) );
  HA1_R03C09 : ha port map (Cout=>HA1_R03C09_C, Sum=>HA1_R03C09_S, A=>PP3(3), B=>PP4(1) );

  FA1_R00C08 : fa port map (Cout=>FA1_R00C08_C, Sum=>FA1_R00C08_S, A=>PP0(8), B=>PP1(6), C=>PP2(4) );
  FA1_R03C08 : fa port map (Cout=>FA1_R03C08_C, Sum=>FA1_R03C08_S, A=>PP3(2), B=>PP4(0), C=>booth_negtive(4) );

  FA1_R00C07 : fa port map (Cout=>FA1_R00C07_C, Sum=>FA1_R00C07_S, A=>PP0(7), B=>PP1(5), C=>PP2(3) );
  FA1_R00C06 : fa port map (Cout=>FA1_R00C06_C, Sum=>FA1_R00C06_S, A=>PP0(6), B=>PP1(4), C=>PP2(2) );
  HA1_R03C06 : ha port map (Cout=>HA1_R03C06_C, Sum=>HA1_R03C06_S, A=>PP3(0), B=>booth_negtive(3) );

  FA1_R00C05 : fa port map (Cout=>FA1_R00C05_C, Sum=>FA1_R00C05_S, A=>PP0(5), B=>PP1(3), C=>PP2(1) );
  FA1_R00C04 : fa port map (Cout=>FA1_R00C04_C, Sum=>FA1_R00C04_S, A=>PP0(4), B=>PP1(2), C=>PP2(0) );

  FA1_R00C02 : fa port map (Cout=>FA1_R00C02_C, Sum=>FA1_R00C02_S, A=>PP0(2), B=>PP1(0), C=>booth_negtive(1) );

  --WCSA step#2

  FA2_R00C15 : fa port map (Cout=>FA2_R00C15_C, Sum=>FA2_R00C15_S, A=>pp_sign_3_not, B=>PP4(7), C=>FA1_R00C14_C );

  HA2_R00C14 : ha port map (Cout=>HA2_R00C14_C, Sum=>HA2_R00C14_S, A=>FA1_R00C14_S, B=>FA1_R00C13_C );
  HA2_R00C13 : ha port map (Cout=>HA2_R00C13_C, Sum=>HA2_R00C13_S, A=>FA1_R00C13_S, B=>FA1_R00C12_C );

  FA2_R00C12 : fa port map (Cout=>FA2_R00C12_C, Sum=>FA2_R00C12_S, A=>FA1_R00C12_S, B=>FA1_R00C11_C, C=> HA1_R03C11_C );
  FA2_R00C11 : fa port map (Cout=>FA2_R00C11_C, Sum=>FA2_R00C11_S, A=>FA1_R00C11_S, B=>FA1_R00C10_C, C=> HA1_R03C11_S );
  FA2_R00C10 : fa port map (Cout=>FA2_R00C10_C, Sum=>FA2_R00C10_S, A=>FA1_R00C10_S, B=>FA1_R00C09_C, C=> HA1_R03C10_S );
  FA2_R00C09 : fa port map (Cout=>FA2_R00C09_C, Sum=>FA2_R00C09_S, A=>FA1_R00C09_S, B=>FA1_R00C08_C, C=> HA1_R03C09_S );
  FA2_R00C08 : fa port map (Cout=>FA2_R00C08_C, Sum=>FA2_R00C08_S, A=>FA1_R00C08_S, B=>FA1_R00C07_C, C=> FA1_R03C08_S );
  FA2_R00C07 : fa port map (Cout=>FA2_R00C07_C, Sum=>FA2_R00C07_S, A=>FA1_R00C07_S, B=>FA1_R00C06_C, C=> HA1_R03C06_C );
  FA2_R00C06 : fa port map (Cout=>FA2_R00C06_C, Sum=>FA2_R00C06_S, A=>FA1_R00C06_S, B=>FA1_R00C05_C, C=> HA1_R03C06_S );

  FA2_R00C03 : fa port map (Cout=> FA2_R00C03_C , Sum=> FA2_R00C03_S , A=>PP0(3) , B=>PP1(1) , C=>FA1_R00C02_C );

  -- WCSA step#3
  HA3_R00C15 : ha port map (Cout=> HA3_R00C15_C , Sum=> HA3_R00C15_S , A=> FA2_R00C15_S , B=> HA2_R00C14_C );
  HA3_R00C14 : ha port map (Cout=> HA3_R00C14_C , Sum=> HA3_R00C14_S , A=> HA2_R00C14_S , B=> HA2_R00C13_C );
  HA3_R00C13 : ha port map (Cout=> HA3_R00C13_C , Sum=> HA3_R00C13_S , A=> HA2_R00C13_S , B=> FA2_R00C12_C );
  FA3_R00C12 : fa port map (Cout=> FA3_R00C12_C , Sum=> FA3_R00C12_S , A=> FA2_R00C12_S , B=> FA2_R00C11_C , C=> PP4(4) );
  FA3_R00C11 : fa port map (Cout=> FA3_R00C11_C , Sum=> FA3_R00C11_S , A=> FA2_R00C11_S , B=> FA2_R00C10_C , C=> HA1_R03C10_C );
  FA3_R00C10 : fa port map (Cout=> FA3_R00C10_C , Sum=> FA3_R00C10_S , A=> FA2_R00C10_S , B=> FA2_R00C09_C , C=> HA1_R03C09_C );
  FA3_R00C09 : fa port map (Cout=> FA3_R00C09_C , Sum=> FA3_R00C09_S , A=> FA2_R00C09_S , B=> FA2_R00C08_C , C=> FA1_R03C08_C );

  HA3_R00C08 : ha port map (Cout=> HA3_R00C08_C , Sum=> HA3_R00C08_S , A=> FA2_R00C08_S , B=> FA2_R00C07_C );
  FA3_R00C07 : fa port map (Cout=> FA3_R00C07_C , Sum=> FA3_R00C07_S , A=> FA2_R00C07_S , B=> FA2_R00C06_C , C=> PP3(1) );

  HA3_R00C05 : ha port map (Cout=> HA3_R00C05_C , Sum=> HA3_R00C05_S , A=> FA1_R00C05_S , B=> FA1_R00C04_C );
  FA3_R00C04 : fa port map (Cout=> FA3_R00C04_C , Sum=> FA3_R00C04_S , A=> FA1_R00C04_S , B=> booth_negtive(2) , C=>FA2_R00C03_C );

  csa_a(0) <= PP0(0);
  csa_b(0) <= booth_negtive(0);
  csa_a(1) <= PP0(1);
  csa_b(1) <= '0';
  csa_a(2) <= FA1_R00C02_S;
  csa_b(2) <= '0';
  csa_a(3) <= FA2_R00C03_S;
  csa_b(3) <= '0';
 
  csa_a(4) <= FA3_R00C04_S;
  csa_b(4) <= '0';
 
  csa_a(5) <= HA3_R00C05_S;
  csa_b(5) <= FA3_R00C04_C;
  csa_a(6) <= FA2_R00C06_S;
  csa_b(6) <= HA3_R00C05_C;
  csa_a(7) <= FA3_R00C07_S;
  csa_b(7) <= '0';
  csa_a(8) <= HA3_R00C08_S;
  csa_b(8) <= FA3_R00C07_C;
  csa_a(9) <= FA3_R00C09_S;
  csa_b(9) <= HA3_R00C08_C;
  csa_a(10) <= FA3_R00C10_S;
  csa_b(10) <= FA3_R00C09_C;
  csa_a(11) <= FA3_R00C11_S;
  csa_b(11) <= FA3_R00C10_C;
  csa_a(12) <= FA3_R00C12_S;
  csa_b(12) <= FA3_R00C11_C;
  csa_a(13) <= HA3_R00C13_S;
  csa_b(13) <= FA3_R00C12_C;
  csa_a(14) <= HA3_R00C14_S;
  csa_b(14) <= HA3_R00C13_C;
  csa_a(15) <= HA3_R00C15_S;
  csa_b(15) <= HA3_R00C14_C;

end MPY8x8_ARCH; 



---------------------------------------------------------------------------
----			MPY16x16 	 	  			---	
---------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;


entity MPY16X16 is 
	port (
		clk		: in	std_logic;  
		IHRST		: in	std_logic; 
		ILRST		: in	std_logic;
		FSEL		: in	std_logic; 
		GSEL		: in 	std_logic;
		HSEL		: in 	std_logic; 
		JKSEL		: in   	std_logic;
		MPY_8X8_MODE	: in   	std_logic;
		ASGND		: in   	std_logic;
		BSGND 		: in   	std_logic;
		A		: in   	std_logic_vector ( 15 downto 0);
		B		: in   	std_logic_vector ( 15 downto 0);
		OH_8X8		: out	std_logic_vector ( 15 downto 0);
		OL_8X8		: out 	std_logic_vector ( 15 downto 0);
		O_16X16		: out   std_logic_vector ( 31 downto 0)
	);
end MPY16X16;  

architecture MPY16X16_ARCH of MPY16X16 is 

 component MPY8x8 is 
	port 	(
		csa_a		: out std_logic_vector( 15 downto 0); 
		csa_b		: out std_logic_vector( 15 downto 0);
		multiplicand    : in  std_logic_vector( 7 downto 0);
		multiplier      : in  std_logic_vector( 7 downto 0); 
		signed_MPD      : std_logic ;    
		signed_MPR      : std_logic
		);
 end component;

 
 component  fcla16 is
        port  (
                Sum     : out   std_logic_vector( 15 downto 0);
                G       : out   std_logic ;
                P       : out   std_logic ;
                A       : in    std_logic_vector( 15 downto 0 );
                B       : in    std_logic_vector( 15 downto 0 );
                Cin     : in    std_logic
                );
 end component; 

 component fcla8 is
        port
          (
                Sum     : out   std_logic_vector( 7 downto 0);
                G       : out   std_logic ;
                P       : out   std_logic ;
                A       : in    std_logic_vector( 7 downto 0);
                B       : in    std_logic_vector( 7 downto 0);
                Cin     : in    std_logic
          );
  end component; 


 component fa is
        port (
                 A      : in    std_logic ;
                 B      : in    std_logic ;
                 C      : in    std_logic ;
                 Sum    : out   std_logic ;
                 Cout   : out   std_logic
               );

 end component; 

  signal  	csa_rega, csa_regb 	: std_logic_vector( 31 downto 0);
  signal  	pp_out		 	: std_logic_vector(152 downto 0);

  signal	MPYG_mpd, MPYG_mpr 	: std_logic_vector( 7 downto 0);
  signal	MPYJ_mpd, MPYJ_mpr	: std_logic_vector( 7 downto 0);
  signal	MPYF_mpd, MPYF_mpr	: std_logic_vector( 7 downto 0);
  signal	MPYK_mpd, MPYK_mpr      : std_logic_vector( 7 downto 0);
  signal	MPYG_MPD_sign, MPYG_MPR_sign : std_logic ;
  signal	MPYJ_MPD_sign, MPYJ_MPR_sign : std_logic ;
  signal	MPYF_MPD_sign, MPYF_MPR_sign : std_logic ;
  signal	MPYK_MPD_sign, MPYK_MPR_sign : std_logic ;

  signal	MPYG_csa_a, MPYG_csa_b : std_logic_vector(15 downto 0);
  signal	MPYJ_csa_a, MPYJ_csa_b : std_logic_vector(15 downto 0);
  signal	MPYF_csa_a, MPYF_csa_b : std_logic_vector(15 downto 0);
  signal	MPYK_csa_a, MPYK_csa_b : std_logic_vector(15 downto 0) ;
  signal	MPYG_o, MPYG_out : std_logic_vector(15 downto 0) ;
  signal	MPYJ_o, MPYJ_out : std_logic_vector(15 downto 0) ;
  signal	MPYF_o, MPYF_out : std_logic_vector(15 downto 0) ;
  signal	MPYK_o, MPYK_out : std_logic_vector(15 downto 0);
  signal	MPYG_oreg, MPYJ_oreg : std_logic_vector(15 downto 0);
  signal	MPYF_oreg, MPYK_oreg : std_logic_vector(15 downto 0);
  signal	MPYJ_out_sign, MPYK_out_sign : std_logic ;
  signal	MPYJK_g, MPYJK_p : std_logic ;


  signal 	MPYG_cla_ina, MPYG_cla_inb : std_logic_vector(15 downto 0) ;
  signal 	CLA16_G_g, CLA16_G_p, MPYG_ci : std_logic ;
  signal        dangle_g_nodeJ, dangle_p_nodeJ : std_logic ; 
  signal 	dangle_g_nodeF, dangle_p_nodeF : std_logic ; 
  signal 	dangle_g_nodeK, dangle_p_nodeK: std_logic ; 

  signal  	csa_oc : std_logic_vector(23 downto 0) ;
  signal 	csa_os : std_logic_vector(23 downto 0) ;
  signal  	MPYJK_g_b : std_logic ;


 signal  	mpy16_reg : std_logic_vector(31 downto 0);


  signal 	cla_ina : std_logic_vector(23 downto 0) ;
  signal 	cla_inb : std_logic_vector(23 downto 0) ;
  signal        cla_o : std_logic_vector(23 downto 0) ;
  signal 	cla24_g0, cla24_p0 : std_logic ;
  signal        cla24_g1, cla24_p1 : std_logic ;
  signal        cla24_cin, cla24_16_cout : std_logic ;

begin 
 --
  MPYG_mpd <= A(7 downto 0);
  MPYG_mpr <= B(7 downto 0);
  process (MPY_8X8_MODE, ASGND) 
   begin 		
	case (MPY_8X8_MODE) is 
	when '0' => MPYG_MPD_sign <= '0'; 	
	when '1' => MPYG_MPD_sign <= ASGND ; 
	when others => MPYG_MPD_sign <= '0'; 
	end case; 
   end process ; 	

  process (MPY_8X8_MODE, BSGND) 
   begin 		
	case (MPY_8X8_MODE) is 
	when '0' => MPYG_MPR_sign <= '0'; 	
	when '1' => MPYG_MPR_sign <= BSGND ; 
	when others => MPYG_MPR_sign <= '0'; 
	end case; 
   end process ;	

   MPYJ_mpd <= A(7 downto 0);
   MPYJ_mpr <= B(15 downto 8);
   MPYJ_MPD_sign <= '0';
   MPYJ_MPR_sign <= BSGND;
   --
   MPYF_mpd <= A(15 downto 8);
   MPYF_mpr <= B(15 downto 8);
   MPYF_MPD_sign <= ASGND;
   MPYF_MPR_sign <= BSGND;
   --
  MPYK_mpd <= A(15 downto 8);
  MPYK_mpr <= B(7 downto 0);
  MPYK_MPD_sign <= ASGND;
  MPYK_MPR_sign <= '0'; 
  --
   process(BSGND, MPYJ_out(15) ) 
   begin
    case (BSGND) is 	
	when '0' => MPYJ_out_sign <= '0';  
        when '1' =>  MPYJ_out_sign <= MPYJ_out(15); 
	when others => MPYJ_out_sign <= '0';  
    end case; 	
   end process; 		


   process(ASGND, MPYK_out(15) ) 
   begin
    case (ASGND) is 	
	when '0' => MPYK_out_sign <= '0';  
        when '1' =>  MPYK_out_sign <= MPYK_out(15); 
	when others => MPYK_out_sign <= '0';  
    end case; 	
   end process; 		

  --
  MPYJK_g <= MPYJ_out_sign and MPYK_out_sign;
  MPYJK_p <= MPYJ_out_sign xor MPYK_out_sign;
  --
 MPY_G: MPY8x8 port map (csa_a=> MPYG_csa_a ,csa_b=> MPYG_csa_b ,multiplicand=> MPYG_mpd ,multiplier=> MPYG_mpr ,signed_MPD=> MPYG_MPD_sign ,signed_MPR=> MPYG_MPR_sign );
 MPY_J: MPY8x8 port map ( csa_a=> MPYJ_csa_a ,csa_b=> MPYJ_csa_b ,multiplicand=> MPYJ_mpd ,multiplier=> MPYJ_mpr ,signed_MPD=> MPYJ_MPD_sign ,signed_MPR=> MPYJ_MPR_sign );
 MPY_F: MPY8x8 port map (csa_a=> MPYF_csa_a ,csa_b=> MPYF_csa_b ,multiplicand=> MPYF_mpd ,multiplier=> MPYF_mpr ,signed_MPD=> MPYF_MPD_sign ,signed_MPR=>MPYF_MPR_sign );
 MPY_K: MPY8x8 port map (csa_a=> MPYK_csa_a ,csa_b=> MPYK_csa_b ,multiplicand=> MPYK_mpd ,multiplier=> MPYK_mpr ,signed_MPD=> MPYK_MPD_sign ,signed_MPR=>MPYK_MPR_sign );


  MPYG_cla_ina <= MPYG_csa_a;
  MPYG_cla_inb <= MPYG_csa_b;

  MPYG_ci <= '0';

  CLA16_G: fcla16  port map 
  (
  	Sum=> MPYG_o(15 downto 0) ,
  	A=> MPYG_cla_ina(15 downto 0) ,
  	B=> MPYG_cla_inb(15 downto 0) , 
  	G=> CLA16_G_g,
  	P=> CLA16_G_p,
  	Cin=>MPYG_ci
  );
  
  CLA16_J: fcla16 port map (
  	Sum=> MPYJ_o(15 downto 0),
  	A=> MPYJ_csa_a(15 downto 0),
  	B=> MPYJ_csa_b(15 downto 0), 
  	Cin=>'0',
  	G=>dangle_g_nodeJ,
  	P=>dangle_p_nodeJ
  );
  
  
  
  CLA16_F : fcla16  port map (
  	Sum=>MPYF_o(15 downto 0) ,
  	A=> MPYF_csa_a(15 downto 0),
  	B=> MPYF_csa_b(15 downto 0) , 
  	Cin=>'0',
  	G=>dangle_g_nodeF,
  	P=>dangle_p_nodeF
  );
  
  
  CLA16_K : fcla16 port map(
  Sum=>MPYK_o(15 downto 0) ,
  A=> MPYK_csa_a(15 downto 0) ,
  B=> MPYK_csa_b(15 downto 0) , 
  Cin=> '0',
  G=>dangle_g_nodeK, 
  P=>dangle_p_nodeK
  );
  

  process(clk,IHRST) 
  begin 
	if(IHRST='1') then 
		MPYF_oreg <= (others => '0'); 
	elsif rising_edge(clk) then 
		MPYF_oreg <= MPYF_o; 
	end if ;
  end process; 

  process(clk,MPY_8X8_MODE,IHRST) 
  begin 
	if(IHRST='1') then 
		MPYJ_oreg <= (others => '0'); 
	elsif (MPY_8X8_MODE ='1') then 
		MPYJ_oreg <=  MPYJ_oreg;  
	elsif rising_edge(clk) then 
		MPYJ_oreg <= MPYJ_o; 
	end if ;
  end process; 

  process(clk,MPY_8X8_MODE,ILRST) 
  begin 
	if(ILRST='1') then 
		MPYK_oreg <= (others => '0'); 
	elsif (MPY_8X8_MODE ='1') then 
		MPYK_oreg <=  MPYK_oreg;  
	elsif rising_edge(clk) then 
		MPYK_oreg <= MPYK_o; 
	end if ;
  end process; 

 
  process(clk,ILRST) 
  begin 
	if(ILRST='1') then 
		MPYG_oreg <= (others => '0'); 
	elsif rising_edge(clk) then 
		MPYG_oreg <= MPYG_o; 
	end if ;
  end process; 

  
   process(GSEL, MPYG_oreg, MPYG_o ) 
   begin
    case (GSEL) is 	
	when '0' => MPYG_out <= MPYG_o ;  
        when '1' =>  MPYG_out <= MPYG_oreg ; 
	when others => MPYG_out <= (others => '0');  
    end case; 	
   end process; 	


   process(JKSEL, MPYJ_oreg, MPYJ_o ) 
   begin
    case (JKSEL) is 	
	when '0' => MPYJ_out <= MPYJ_o ;  
        when '1' =>  MPYJ_out <= MPYJ_oreg ; 
	when others => MPYJ_out <= (others => '0');  
    end case; 	
   end process; 	


   process(JKSEL, MPYF_oreg, MPYF_o ) 
   begin
    case (JKSEL) is 	
	when '0' => MPYF_out <= MPYF_o ;  
        when '1' =>  MPYF_out <= MPYF_oreg ; 
	when others => MPYF_out <= (others => '0');  
    end case; 	
   end process; 	


   process(FSEL, MPYK_oreg, MPYK_o ) 
   begin
    case (FSEL) is 	
	when '0' => MPYK_out <= MPYK_o ;  
        when '1' =>  MPYK_out <= MPYK_oreg ; 
	when others => MPYK_out <= (others => '0');  
    end case; 	
   end process; 	
  	
   MPYJK_g_b <= not(MPYJK_g);

  csa_os(23) <= MPYJK_p xor  MPYF_out(15);
  csa_oc(23) <= not(MPYJK_g_b and not(MPYJK_p and MPYF_out(15)));
  csa_os(22) <= MPYJK_p xor MPYF_out(14);
  csa_oc(22) <= not(MPYJK_g_b and not(MPYJK_p and MPYF_out(14)));
  csa_os(21) <= MPYJK_p xor MPYF_out(13);
  csa_oc(21) <= not(MPYJK_g_b and  not(MPYJK_p and  MPYF_out(13)));
  csa_os(20) <= MPYJK_p xor MPYF_out(12);
  csa_oc(20) <= not(MPYJK_g_b and not(MPYJK_p and MPYF_out(12)));
  csa_os(19) <= MPYJK_p xor MPYF_out(11);
  csa_oc(19) <= not(MPYJK_g_b and  not(MPYJK_p and MPYF_out(11)));
  csa_os(18) <= MPYJK_p xor MPYF_out(10);
  csa_oc(18) <= not(MPYJK_g_b and not(MPYJK_p and MPYF_out(10)));
  csa_os(17) <= MPYJK_p xor MPYF_out(9);
  csa_oc(17) <= not(MPYJK_g_b and not(MPYJK_p and MPYF_out(9)));
  csa_os(16) <= MPYJK_p xor MPYF_out(8);
  csa_oc(16) <= not(MPYJK_g_b and  not(MPYJK_p and MPYF_out(8)));

  FA1_R00C15: fa port map (Cout=>csa_oc(15), Sum=>csa_os(15), A=> MPYJ_out(15) , B=>MPYK_out(15) , C=>MPYF_out(7) );
  FA1_R00C14: fa port map (Cout=>csa_oc(14), Sum=>csa_os(14), A=> MPYJ_out(14) , B=>MPYK_out(14) , C=>MPYF_out(6) );
  FA1_R00C13: fa port map (Cout=>csa_oc(13), Sum=>csa_os(13), A=> MPYJ_out(13) , B=>MPYK_out(13) , C=>MPYF_out(5) );
  FA1_R00C12: fa port map (Cout=>csa_oc(12), Sum=>csa_os(12), A=> MPYJ_out(12) , B=>MPYK_out(12) , C=>MPYF_out(4) );
  FA1_R00C11: fa port map (Cout=>csa_oc(11), Sum=>csa_os(11), A=> MPYJ_out(11) , B=>MPYK_out(11) , C=>MPYF_out(3) );
  FA1_R00C10: fa port map (Cout=>csa_oc(10), Sum=>csa_os(10), A=> MPYJ_out(10) , B=>MPYK_out(10) , C=>MPYF_out(2) );
  FA1_R00C09: fa port map (Cout=>csa_oc(9),  Sum=>csa_os(9),  A=> MPYJ_out(9) ,  B=>MPYK_out(9) ,  C=>MPYF_out(1) );
  FA1_R00C08: fa port map (Cout=>csa_oc(8),  Sum=>csa_os(8),  A=> MPYJ_out(8) ,  B=>MPYK_out(8) ,  C=>MPYF_out(0) );

  FA1_R00C07: fa port map (Cout=>csa_oc(7), Sum=>csa_os(7), A=> MPYG_out(15) , B=>MPYJ_out(7) , C=> MPYK_out(7) );
  FA1_R00C06: fa port map (Cout=>csa_oc(6), Sum=>csa_os(6), A=> MPYG_out(14) , B=>MPYJ_out(6) , C=> MPYK_out(6) );
  FA1_R00C05: fa port map (Cout=>csa_oc(5), Sum=>csa_os(5), A=> MPYG_out(13) , B=>MPYJ_out(5) , C=> MPYK_out(5) );
  FA1_R00C04: fa port map (Cout=>csa_oc(4), Sum=>csa_os(4), A=> MPYG_out(12) , B=>MPYJ_out(4) , C=> MPYK_out(4) );
  FA1_R00C03: fa port map (Cout=>csa_oc(3), Sum=>csa_os(3), A=> MPYG_out(11) , B=>MPYJ_out(3) , C=> MPYK_out(3) );
  FA1_R00C02: fa port map (Cout=>csa_oc(2), Sum=>csa_os(2), A=> MPYG_out(10) , B=>MPYJ_out(2) , C=> MPYK_out(2) );
  FA1_R00C01: fa port map (Cout=>csa_oc(1), Sum=>csa_os(1), A=> MPYG_out(9) ,  B=>MPYJ_out(1) , C=> MPYK_out(1) );
  FA1_R00C00: fa port map (Cout=>csa_oc(0), Sum=>csa_os(0), A=> MPYG_out(8) ,  B=>MPYJ_out(0) , C=> MPYK_out(0) );


 cla_ina <= csa_os;
 cla_inb <= csa_oc(22 downto 0) & '0';
 cla24_cin <= '0';

 CLA24_16 : fcla16  port map (
  	Sum=> cla_o(15 downto 0),
  	G=>	cla24_g0,
  	P=>cla24_p0, 
  	A=>cla_ina(15 downto 0),
  	B=>cla_inb(15 downto 0), 
  	Cin=>cla24_cin
 );

 cla24_16_cout <= not(not(cla24_g0) and not(cla24_p0 and cla24_cin));

 CLA24_8 :  fcla8  port map (
   Sum=>	cla_o(23 downto 16),
   G => 	cla24_g1,
   P => 	cla24_p1, 
   A => 	cla_ina(23 downto 16),
   B => 	cla_inb(23 downto 16), 
   Cin => 	cla24_16_cout
 );

--

  process(clk,ILRST,MPY_8x8_MODE) 
  begin 
	if(ILRST='1') then 
		mpy16_reg  <= (others => '0'); 
	elsif rising_edge(clk) then 
		if(MPY_8X8_MODE = '1') then 
		        mpy16_reg <= mpy16_reg ; 
		else 
			mpy16_reg <= cla_o & MPYG_out(7 downto 0);
		end if ;	
		
	end if ;
  end process; 

--
  process(HSEL, mpy16_reg , cla_o,MPYG_out) 
  begin 
	case (HSEL) is 
	when '0' => O_16X16 <= cla_o & MPYG_out(7 downto 0); 
	when '1' => O_16X16 <= mpy16_reg ; 
	when others =>  O_16X16 <= (others => '0'); 
	end case; 
  end process;
 
	
--
   OH_8X8 <= MPYF_out(15 downto 0);
   OL_8X8 <= MPYG_out(15 downto 0);
--
end MPY16X16_ARCH; 

---------------------------------------------------------
-----------     mac16_physical					   ------
---------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;


entity  mac16_physical  is 
	port  (
	 	CLK				: in	std_logic ; 
	 	IHRST				: in	std_logic ;
	 	ILRST				: in	std_logic ;
	 	OHRST				: in	std_logic ;
	 	OLRST				: in	std_logic ;
	 	A 				: in	std_logic_vector (15 downto 0);
	 	B 				: in	std_logic_vector (15 downto 0);
	 	C 				: in	std_logic_vector (15 downto 0);
	 	D 				: in	std_logic_vector (15 downto 0);
	    	CBIT				: in	std_logic_vector (24 downto 0);
	    	AHLD				: in	std_logic ;
	 	BHLD				: in	std_logic ;
	 	CHLD				: in	std_logic ;
	 	DHLD				: in	std_logic ;
	 	OHHLD				: in	std_logic ;
	 	OLHLD				: in	std_logic ;
		OHADS				: in	std_logic ;
	 	OLADS				: in	std_logic ;
	 	OHLDA				: in	std_logic ;
	 	OLLDA				: in	std_logic ;
	 	CICAS				: in	std_logic ;
	 	CI				: in	std_logic ;
	 	SIGNEXTIN			: in	std_logic ;
	 	SIGNEXTOUT			: out	std_logic ;
	 	COCAS				: out	std_logic ;
	 	CO				: out 	std_logic ;
	 	O				: out	std_logic_vector (31 downto 0)	
    );
end mac16_physical; 
	

architecture mac16_physical_arch of mac16_physical is  

	component REG_BYPASS_MUX is 
  	generic ( 
		DATA_WIDTH : integer 		 := 16 ) ; 
	port 	(
		CLK	   : in std_logic ; 
		RST 	   : in std_logic; 
		ENA	   : in std_logic ;
		D	   : in  std_logic_vector(DATA_WIDTH-1 downto 0);
		SELM	   : in std_logic ;
		Q          : out  std_logic_vector(DATA_WIDTH-1	downto 0)  
		); 
	end component; 	 


	component  MULT_ACCUM is 
	port  (
		DIRECT_INPUT	: in std_logic_vector ( 15 downto 0); 
		MULT_INPUT	: in std_logic_vector ( 15 downto 0);
    		MULT_8x8	: in std_logic_vector ( 15 downto 0);	
		MULT_16x16	: in std_logic_vector ( 15 downto 0);
		ADDSUB		: in std_logic ; 
		CLK		: in std_logic ;
    		CICAS		: in std_logic ;
    		CI		: in std_logic ;
		SIGNEXTIN	: in std_logic ;
		SIGNEXTOUT	: out std_logic ;
    		LDA		: in std_logic ; 
    		RST		: in std_logic ;
    		ENA		: in std_logic ;
    		COCAS		: out std_logic ;
    		CO		: out std_logic ;
    		O		: out std_logic_vector ( 15 downto 0);
		OUTMUX_SEL	: in std_logic_vector ( 1 downto 0);
		CARRYMUX_SEL	: in std_logic_vector ( 1 downto 0);
		ADDER_A_IN_SEL  : in std_logic;
		ADDER_B_IN_SEL  : in std_logic_vector ( 1 downto 0)
    		);
	end component; 

	component MPY16X16 is 
	port (
		clk		: in	std_logic;  
		IHRST		: in	std_logic; 
		ILRST		: in	std_logic;
		FSEL		: in	std_logic; 
		GSEL		: in 	std_logic;
		HSEL		: in 	std_logic; 
		JKSEL		: in   	std_logic;
		MPY_8X8_MODE	: in   	std_logic;
		ASGND		: in   	std_logic;
		BSGND 		: in   	std_logic;
		A		: in   	std_logic_vector ( 15 downto 0);
		B		: in   	std_logic_vector ( 15 downto 0);
		OH_8X8		: out	std_logic_vector ( 15 downto 0);
		OL_8X8		: out 	std_logic_vector ( 15 downto 0);
		O_16X16		: out   std_logic_vector ( 31 downto 0)
	);
	end component;  


	signal AENA, BENA, CENA, DENA, OHENA, OLENA 			: std_logic ;
	signal ASEL, BSEL, CSEL, DSEL, FSEL, JKSEL, GSEL, HSEL 		: std_logic ;
	signal OHADDA_SEL, OLADDA_SEL, MPY_8X8_MODE, ASGND, BSGND 	: std_logic ;
	signal OHOMUX_SEL, OLOMUX_SEL, OHADDB_SEL, OLADDB_SEL, OHCARRYMUX_SEL, OLCARRYMUX_SEL : std_logic_vector( 1 downto 0 );

	signal  REG_A 	: std_logic_vector( 15 downto 0);
	signal  REG_B 	: std_logic_vector( 15 downto 0);
	signal  REG_C 	: std_logic_vector( 15 downto 0);
	signal  REG_D 	: std_logic_vector( 15 downto 0);

	signal  OH_8X8	: std_logic_vector ( 15 downto 0);
	signal  OL_8X8	: std_logic_vector ( 15 downto 0);
	signal  O_16X16	: std_logic_vector ( 31 downto 0);

	signal MAC16_SIGNOUT_L, MAC16_SIGNOUT_H		: std_logic ;  
	signal COCAS_L , CO_L 				: std_logic ;

begin 

	 AENA <= not(AHLD);
	 BENA <= not(BHLD);
	 CENA <= not(CHLD);
	 DENA  <= not(DHLD);
	 OHENA <= not(OHHLD);
	 OLENA <= not(OLHLD);
	 ASEL <= CBIT(1);
	 BSEL <= CBIT(2);
	 CSEL <= CBIT(0);
	 DSEL <= CBIT(3);
	 FSEL <= CBIT(4);
	 JKSEL <= CBIT(6);
	 GSEL <= CBIT(5);
	 HSEL <= CBIT(7);
	OHOMUX_SEL(1 downto 0) <= CBIT(9 downto 8);	
	OLOMUX_SEL(1 downto 0) <= CBIT(16 downto 15);	
	OHADDA_SEL <= CBIT(12);
	OLADDA_SEL <= CBIT(19);
	OHADDB_SEL(1 downto 0) <= CBIT(11 downto 10) ;	
	OLADDB_SEL(1 downto 0)  <= CBIT(18 downto 17) ;	
	OHCARRYMUX_SEL(1 downto 0) <= CBIT(14 downto 13);
	OLCARRYMUX_SEL(1 downto 0) <= CBIT(21 downto 20);
	MPY_8X8_MODE <= CBIT(22);
	ASGND <= CBIT(23);
	BSGND <= CBIT(24);

	
	SIGNEXTOUT <= MAC16_SIGNOUT_H;

A_REG : REG_BYPASS_MUX  port map  (
	D    		=> A ,
	Q    		=> REG_A ,
	ENA  		=> AENA ,
	CLK  		=> CLK,
	RST  		=> IHRST,
	SELM 		=> ASEL 
	); 

B_REG : REG_BYPASS_MUX  port map  (
	 D		=>  B ,
	 Q		=>  REG_B ,
	 ENA 		=> BENA ,
	 CLK 		=> CLK ,
	 RST 		=> ILRST ,
	 SELM 		=> BSEL 
	); 

C_REG : REG_BYPASS_MUX port map   (
	 D 		=> C,
	 Q 		=> REG_C,
	 ENA 		=> CENA ,
	 CLK 		=> CLK ,
	 RST 		=> IHRST ,
	SELM 		=> CSEL 
	); 

D_REG : REG_BYPASS_MUX  port map (
	 D		=> D ,
	 Q		=> REG_D,
	 ENA 		=> DENA ,
	 CLK 		=> CLK ,
	 RST 		=> ILRST,
	 SELM 		=> DSEL  
	); 

HI_MAC : MULT_ACCUM  port map  (
	DIRECT_INPUT 		=> REG_C,
	MULT_INPUT 		=> REG_A,
	MULT_8x8 		=> OH_8X8(15 downto 0),
	MULT_16x16 		=> O_16X16(31 downto 16),
	ADDSUB 			=> OHADS,
	CLK 			=> CLK,
	CICAS 			=> COCAS_L,
	CI 			=> CO_L,
	SIGNEXTIN 		=> MAC16_SIGNOUT_L ,
	SIGNEXTOUT 		=> MAC16_SIGNOUT_H ,
	LDA 			=> OHLDA,
	RST 			=> OHRST,
	ENA 			=> OHENA,
	COCAS 			=> COCAS,
	CO 			=> CO,
	O 			=> O(31 downto 16),
	OUTMUX_SEL 		=> OHOMUX_SEL(1 downto 0),
	ADDER_A_IN_SEL 		=> OHADDA_SEL,
	ADDER_B_IN_SEL 		=> OHADDB_SEL(1 downto 0),
	CARRYMUX_SEL 		=> OHCARRYMUX_SEL(1 downto 0)
    );

LO_MAC : MULT_ACCUM  port map  (
	DIRECT_INPUT  		=> REG_D,
	MULT_INPUT	  	=> REG_B,
	MULT_8x8	  	=> OL_8X8(15 downto 0),
	MULT_16x16	  	=> O_16X16(15 downto 0),
	ADDSUB	      		=> OLADS,
	CLK		      	=> CLK,
	CICAS	      		=> CICAS,
	CI		      	=> CI,
	SIGNEXTIN	  	=> SIGNEXTIN,
	SIGNEXTOUT	  	=> MAC16_SIGNOUT_L,
	LDA			=> OLLDA,
	RST			=> OLRST,
	ENA			=> OLENA,
	COCAS		  	=> COCAS_L,
	CO			=> CO_L,
	O			=> O(15 downto 0),
	OUTMUX_SEL     		=> OLOMUX_SEL(1 downto 0),
	ADDER_A_IN_SEL 		=> OLADDA_SEL,
	ADDER_B_IN_SEL 		=> OLADDB_SEL(1 downto 0),
	CARRYMUX_SEL   		=> OLCARRYMUX_SEL(1 downto 0)
    );
	 
MULTIPLER : MPY16X16  port map  (
	 clk			=> CLK,
	 IHRST			=> IHRST,
	 ILRST			=> ILRST,
	 FSEL			=> FSEL,
	 GSEL			=> GSEL,
	 HSEL			=> HSEL,
	 JKSEL			=> JKSEL,
	 MPY_8X8_MODE		=> MPY_8X8_MODE,
	 ASGND			=> ASGND,
	 BSGND			=> BSGND,
	 A			=> REG_A(15 downto 0),
	 B			=> REG_B(15 downto 0),
	 OH_8X8			=> OH_8X8(15 downto 0),
	 OL_8X8			=> OL_8X8(15 downto 0),
	 O_16X16		=> O_16X16(31 downto 0)
);

end mac16_physical_arch;

---------------------------------------------------------------------------
----			 	SB_MAC16 				---	
---------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use IEEE.numeric_std.all;
--use work.std_logic_SBT.all;


entity SB_MAC16 is
 
	generic ( 	
	
		TimingChecksOn : boolean := true;
		Xon   : boolean := true;
		MsgOn : boolean := true;
		tipd_A		:VitalDelayArrayType01(15 downto 0)  := (others => (0 ns, 0 ns));
		tipd_B		: VitalDelayArrayType01(15 downto 0)  := (others => (0 ns, 0 ns));
		tipd_C		:VitalDelayArrayType01(15 downto 0)  := (others => (0 ns, 0 ns));
		tipd_D		: VitalDelayArrayType01(15 downto 0)  := (others => (0 ns, 0 ns));
		tipd_CLK		: VitalDelayType01 := (0.000 ns, 0.000 ns); 
		tipd_CE		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_IRSTTOP 	: VitalDelayType01 := (0.000 ns, 0.000 ns); 
	    tipd_IRSTBOT 	: VitalDelayType01 := (0.000 ns, 0.000 ns);  
		tipd_ORSTTOP 	: VitalDelayType01 := (0.000 ns, 0.000 ns); 
		tipd_ORSTBOT 	: VitalDelayType01 := (0.000 ns, 0.000 ns); 
		tipd_AHOLD 		:VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_BHOLD		: VitalDelayType01 := (0.000 ns, 0.000 ns); 
		tipd_CHOLD		: VitalDelayType01 := (0.000 ns, 0.000 ns); 
		tipd_DHOLD		: VitalDelayType01 := (0.000 ns, 0.000 ns); 
		tipd_OHOLDTOP	: VitalDelayType01 := (0.000 ns, 0.000 ns); 
		tipd_OHOLDBOT	: VitalDelayType01 := (0.000 ns, 0.000 ns); 
		tipd_OLOADTOP	:VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OLOADBOT	: VitalDelayType01 := (0.000 ns, 0.000 ns); 
		tipd_ADDSUBTOP	: VitalDelayType01 := (0.000 ns, 0.000 ns); 
		tipd_ADDSUBBOT	: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CI		: VitalDelayType01 := (0.000 ns, 0.000 ns); 
		tipd_ACCUMCI		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_SIGNEXTIN	: VitalDelayType01 := (0.000 ns, 0.000 ns);	
		
		tpd_IRSTBOT_O : VitalDelayArrayType01(31 downto 0) := (others => (0.0 ns, 0.0 ns));
		tpd_CLK_O_posedge : VitalDelayArrayType01(31 downto 0) := (others => (0.0 ns, 0.0 ns));
		tpd_ORSTBOT_O : VitalDelayArrayType01(31 downto 0) := (others => (0.0 ns, 0.0 ns));
		tpd_ORSTTOP_O : VitalDelayArrayType01(31 downto 0) := (others => (0.0 ns, 0.0 ns));	
		tpd_CI_O : VitalDelayArrayType01(31 downto 0) := (others => (0.0 ns, 0.0 ns));
		tpd_ADDSUBTOP_O : VitalDelayArrayType01(31 downto 0) := (others => (0.0 ns, 0.0 ns));
		tpd_ADDSUBBOT_O : VitalDelayArrayType01(31 downto 0) := (others => (0.0 ns, 0.0 ns));
		tpd_OLOADTOP_O : VitalDelayArrayType01(31 downto 0) := (others => (0.0 ns, 0.0 ns)); 
		tpd_OLOADBOT_O : VitalDelayArrayType01(31 downto 0) := (others => (0.0 ns, 0.0 ns));
		tpd_A_CO : VitalDelayArrayType01(15 downto 0) := (others => (0.0 ns, 0.0 ns));	
		tpd_A_ACCUMCO : VitalDelayArrayType01(15 downto 0) := (others => (0.0 ns, 0.0 ns));	
		tpd_B_CO : VitalDelayArrayType01(15 downto 0) := (others => (0.0 ns, 0.0 ns));	
		tpd_B_ACCUMCO : VitalDelayArrayType01(15 downto 0) := (others => (0.0 ns, 0.0 ns));	
		tpd_C_CO : VitalDelayArrayType01(15 downto 0) := (others => (0.0 ns, 0.0 ns));	
		tpd_C_ACCUMCO : VitalDelayArrayType01(15 downto 0) := (others => (0.0 ns, 0.0 ns));	
		tpd_D_CO : VitalDelayArrayType01(15 downto 0) := (others => (0.0 ns, 0.0 ns));	
		tpd_D_ACCUMCO : VitalDelayArrayType01(15 downto 0) := (others => (0.0 ns, 0.0 ns));	
		tpd_CI_CO : VitalDelayType01 := (0.000 ns, 0.000 ns);		
		tpd_CI_ACCUMCO : VitalDelayType01 := (0.000 ns, 0.000 ns)	;
		tpd_OLOADTOP_CO : VitalDelayType01 := (0.000 ns, 0.000 ns);		
		tpd_OLOADTOP_ACCUMCO : VitalDelayType01 := (0.000 ns, 0.000 ns);	
		tpd_OLOADBOT_CO : VitalDelayType01 := (0.000 ns, 0.000 ns);		
		tpd_OLOADBOT_ACCUMCO : VitalDelayType01 := (0.000 ns, 0.000 ns)	;	
		tpd_ADDSUBBOT_CO : VitalDelayType01 := (0.000 ns, 0.000 ns);		
		tpd_ADDSUBBOT_ACCUMCO : VitalDelayType01 := (0.000 ns, 0.000 ns)	;	
		tpd_CLK_CO_posedge : VitalDelayType01 := (0.000 ns, 0.000 ns);		
		tpd_CLK_ACCUMCO_posedge : VitalDelayType01 := (0.000 ns, 0.000 ns)	;	
		tpd_ACCUMCI_CO : VitalDelayType01 := (0.000 ns, 0.000 ns);	
		tpd_ACCUMCI_ACCUMCO : VitalDelayType01 := (0.000 ns, 0.000 ns)	;	
		tpd_ACCUMCI_O : VitalDelayArrayType01(31 downto 0) := (others => (0.0 ns, 0.0 ns));
		
		tpd_A_SIGNEXTOUT : VitalDelayArrayType01(15 downto 0) := (others => (0.0 ns, 0.0 ns));
		tpd_B_SIGNEXTOUT : VitalDelayArrayType01(15 downto 0) := (others => (0.0 ns, 0.0 ns));
		tpd_CLK_SIGNEXTOUT_posedge : VitalDelayType01 := (0.000 ns, 0.000 ns);
		tpd_ADDSUBTOP_ACCUMCO                : VitalDelayType01 := (0 ns, 0 ns);
		tpd_ADDSUBTOP_CO                : VitalDelayType01 := (0 ns, 0 ns);
		
		tpd_A_O : VitalDelayArrayType01(511 downto 0):= (others => (0.0 ns, 0.0 ns)); 
		tpd_B_O : VitalDelayArrayType01(511 downto 0) := (others => (0.0 ns, 0.0 ns)); 
		tpd_C_O : VitalDelayArrayType01(511 downto 0) := (others => (0.0 ns, 0.0 ns)); 
		tpd_D_O : VitalDelayArrayType01(511 downto 0) := (others => (0.0 ns, 0.0 ns));

		 tsetup_A_CLK_posedge_posedge : VitalDelayArrayType(15 downto 0)  := (others => 0 ns);
		 tsetup_A_CLK_negedge_posedge : VitalDelayArrayType(15 downto 0)  := (others => 0 ns);
		 tsetup_B_CLK_posedge_posedge : VitalDelayArrayType(15 downto 0)  := (others => 0 ns);
		 tsetup_B_CLK_negedge_posedge : VitalDelayArrayType(15 downto 0)  := (others => 0 ns);
		 tsetup_C_CLK_posedge_posedge : VitalDelayArrayType(15 downto 0)  := (others => 0 ns);
		 tsetup_C_CLK_negedge_posedge : VitalDelayArrayType(15 downto 0)  := (others => 0 ns);
		 tsetup_D_CLK_posedge_posedge : VitalDelayArrayType(15 downto 0)  := (others => 0 ns);
		 tsetup_D_CLK_negedge_posedge : VitalDelayArrayType(15 downto 0)  := (others => 0 ns);		 
		 tsetup_ADDSUBTOP_CLK_posedge_posedge : VitalDelayType := 0 ns;
		 tsetup_ADDSUBTOP_CLK_negedge_posedge : VitalDelayType  := 0 ns;
		 tsetup_ADDSUBBOT_CLK_posedge_posedge : VitalDelayType  := 0 ns;
		 tsetup_ADDSUBBOT_CLK_negedge_posedge : VitalDelayType := 0 ns;
		 tsetup_OLOADTOP_CLK_posedge_posedge : VitalDelayType := 0 ns;
		 tsetup_OLOADTOP_CLK_negedge_posedge : VitalDelayType  := 0 ns;
		 tsetup_OLOADBOT_CLK_posedge_posedge : VitalDelayType  := 0 ns;
		 tsetup_OLOADBOT_CLK_negedge_posedge : VitalDelayType := 0 ns;	
		 tsetup_OHOLDBOT_CLK_posedge_posedge : VitalDelayType := 0 ns;
		 tsetup_OHOLDBOT_CLK_negedge_posedge : VitalDelayType  := 0 ns;
		 tsetup_OHOLDTOP_CLK_posedge_posedge : VitalDelayType  := 0 ns;
		 tsetup_OHOLDTOP_CLK_negedge_posedge : VitalDelayType := 0 ns;	
		 tsetup_AHOLD_CLK_posedge_posedge : VitalDelayType := 0 ns;
		 tsetup_AHOLD_CLK_negedge_posedge : VitalDelayType  := 0 ns;
		 tsetup_BHOLD_CLK_posedge_posedge : VitalDelayType  := 0 ns;
		 tsetup_BHOLD_CLK_negedge_posedge : VitalDelayType := 0 ns;
		 tsetup_CHOLD_CLK_posedge_posedge : VitalDelayType := 0 ns;
		 tsetup_CHOLD_CLK_negedge_posedge : VitalDelayType  := 0 ns;
		 tsetup_DHOLD_CLK_posedge_posedge : VitalDelayType  := 0 ns;
		 tsetup_DHOLD_CLK_negedge_posedge : VitalDelayType := 0 ns;			 
		 tsetup_CI_CLK_posedge_posedge : VitalDelayType  := 0 ns;	  
		 tsetup_CI_CLK_negedge_posedge : VitalDelayType := 0 ns;		 
		 tsetup_ACCUMCI_CLK_posedge_posedge : VitalDelayType  := 0 ns;	  
		 tsetup_ACCUMCI_CLK_negedge_posedge : VitalDelayType := 0 ns;
		
		 thold_A_CLK_posedge_posedge : VitalDelayArrayType(15 downto 0)  := (others => 0 ns);
		 thold_A_CLK_negedge_posedge : VitalDelayArrayType(15 downto 0)  := (others => 0 ns);
		 thold_B_CLK_posedge_posedge : VitalDelayArrayType(15 downto 0)  := (others => 0 ns);
		 thold_B_CLK_negedge_posedge : VitalDelayArrayType(15 downto 0)  := (others => 0 ns);
		 thold_C_CLK_posedge_posedge : VitalDelayArrayType(15 downto 0)  := (others => 0 ns);
		 thold_C_CLK_negedge_posedge : VitalDelayArrayType(15 downto 0)  := (others => 0 ns);
		 thold_D_CLK_posedge_posedge : VitalDelayArrayType(15 downto 0)  := (others => 0 ns);
		 thold_D_CLK_negedge_posedge : VitalDelayArrayType(15 downto 0)  := (others => 0 ns);		 
		 thold_ADDSUBTOP_CLK_posedge_posedge : VitalDelayType := 0 ns;
		 thold_ADDSUBTOP_CLK_negedge_posedge : VitalDelayType  := 0 ns;
		 thold_ADDSUBBOT_CLK_posedge_posedge : VitalDelayType  := 0 ns;
		 thold_ADDSUBBOT_CLK_negedge_posedge : VitalDelayType := 0 ns;
		 thold_OLOADTOP_CLK_posedge_posedge : VitalDelayType := 0 ns;
		 thold_OLOADTOP_CLK_negedge_posedge : VitalDelayType  := 0 ns;
		 thold_OLOADBOT_CLK_posedge_posedge : VitalDelayType  := 0 ns;
		 thold_OLOADBOT_CLK_negedge_posedge : VitalDelayType := 0 ns;
		 thold_OHOLDBOT_CLK_posedge_posedge	: VitalDelayType := 0 ns;
		 thold_OHOLDBOT_CLK_negedge_posedge	: VitalDelayType := 0 ns;  
		  thold_OHOLDTOP_CLK_posedge_posedge	: VitalDelayType := 0 ns;
		  thold_OHOLDTOP_CLK_negedge_posedge	: VitalDelayType := 0 ns;
		 thold_AHOLD_CLK_posedge_posedge : VitalDelayType := 0 ns;
		 thold_AHOLD_CLK_negedge_posedge : VitalDelayType  := 0 ns;
		 thold_BHOLD_CLK_posedge_posedge : VitalDelayType  := 0 ns;
		 thold_BHOLD_CLK_negedge_posedge : VitalDelayType := 0 ns;
		 thold_CHOLD_CLK_posedge_posedge : VitalDelayType := 0 ns;
		 thold_CHOLD_CLK_negedge_posedge : VitalDelayType  := 0 ns;
		 thold_DHOLD_CLK_posedge_posedge : VitalDelayType  := 0 ns;
		 thold_DHOLD_CLK_negedge_posedge : VitalDelayType := 0 ns;			 
		 thold_CI_CLK_posedge_posedge : VitalDelayType  := 0 ns;
		 thold_CI_CLK_negedge_posedge : VitalDelayType := 0 ns;	
		 thold_ACCUMCI_CLK_posedge_posedge : VitalDelayType  := 0 ns;
		 thold_ACCUMCI_CLK_negedge_posedge : VitalDelayType := 0 ns;

		 tpw_CLK_negedge : VitalDelayType := 0 ns;
		 tpw_CLK_posedge : VitalDelayType := 0 ns;
		 tperiod_CLK_posedge : VitalDelayType := 0 ns;


           trecovery_IRSTTOP_CLK_posedge_posedge  : VitalDelayType                   := 0 ns;
           trecovery_IRSTTOP_CLK_negedge_posedge  : VitalDelayType                   := 0 ns;
           tremoval_IRSTTOP_CLK_posedge_posedge   : VitalDelayType                   := 0 ns;
           tremoval_IRSTTOP_CLK_negedge_posedge   : VitalDelayType                   := 0 ns;
           trecovery_IRSTBOT_CLK_posedge_posedge  : VitalDelayType                   := 0 ns;
           trecovery_IRSTBOT_CLK_negedge_posedge  : VitalDelayType                   := 0 ns;
           tremoval_IRSTBOT_CLK_posedge_posedge   : VitalDelayType                   := 0 ns;
           tremoval_IRSTBOT_CLK_negedge_posedge   : VitalDelayType                   := 0 ns;
		   
		   trecovery_ORSTTOP_CLK_posedge_posedge  : VitalDelayType                   := 0 ns;
           trecovery_ORSTTOP_CLK_negedge_posedge  : VitalDelayType                   := 0 ns;
           tremoval_ORSTTOP_CLK_posedge_posedge   : VitalDelayType                   := 0 ns;
           tremoval_ORSTTOP_CLK_negedge_posedge   : VitalDelayType                   := 0 ns;
           trecovery_ORSTBOT_CLK_posedge_posedge  : VitalDelayType                   := 0 ns;
           trecovery_ORSTBOT_CLK_negedge_posedge  : VitalDelayType                   := 0 ns;
           tremoval_ORSTBOT_CLK_posedge_posedge   : VitalDelayType                   := 0 ns;
           tremoval_ORSTBOT_CLK_negedge_posedge   : VitalDelayType                   := 0 ns;
		 
		 
		NEG_TRIGGER 			: bit 		:='0'; 
		 C_REG				: bit 		:='0'; 		-- C0
		 A_REG				: bit 		:='0'; 	    	-- C1 
		 B_REG				: bit 		:='0';		-- C2
		 D_REG 				: bit 		:='0';		-- C3

		 TOP_8x8_MULT_REG		: bit 		:='0'; 	   	-- C4
		 BOT_8x8_MULT_REG		: bit 		:='0';	   	-- C5
		 PIPELINE_16x16_MULT_REG1	: bit 		:='0';		-- C6
		 PIPELINE_16x16_MULT_REG2	: bit 		:='0';		-- C7

		 TOPOUTPUT_SELECT      		: bit_vector(1 downto 0) := "00" ;	-- COMB, ACCUM_REG, MULT_8x8, MULT_16x16 //{C9,C8}   = 00, 01, 10, 11
		 TOPADDSUB_LOWERINPUT  		: bit_vector(1 downto 0) := "00" ; 	-- DATA, MULT_8x8, MULT_16x16, SIGNEXT 	 //{C11,C10} = 00, 01, 10, 11
		 TOPADDSUB_UPPERINPUT  		: bit 			 := '0'  ; 	-- ACCUM_REG, DATAC 		 	 // C12 = 0, 1
		 TOPADDSUB_CARRYSELECT 		: bit_vector(1 downto 0) := "00" ; 	-- LOGIC0,LOGIC1,ACCUMCI,GENERATED_CARRY //{C14, C13} =00, 01, 10, 11

		 BOTOUTPUT_SELECT		: bit_vector(1 downto 0) := "00" ; 	--COMB, ACCUM_REG, MULT_8x8, MULT_16x16  // {C16,C15} =00, 01, 10, 11
		 BOTADDSUB_LOWERINPUT 		: bit_vector(1 downto 0) := "00" ; 	--DATA, MULT_8x8, MULT_16x16, SIGNEXTIN //  {C18,C17} =00, 01, 10, 11
		 BOTADDSUB_UPPERINPUT 		: bit 			 := '0'  ;  	--ACCUM_REG, DATAD   			//  C19 = 0, 1
		 BOTADDSUB_CARRYSELECT 		: bit_vector(1 downto 0) := "00" ; 	--LOGIC0, LOGIC1, ACCUMCI, CI  		//  {C21, C20}=00,01,10,11
		 MODE_8x8 			: bit 			 := '0' ; 	-- C22 

		 A_SIGNED 			: bit 			 := '0' ;  	-- C23
		 B_SIGNED 			: bit 			 := '0'   	-- C24
	);
	port	(

		A		: in 	std_logic_vector(15 downto 0) := x"0000";  
		B		: in    std_logic_vector(15 downto 0) := x"0000"; 	
		C		: in 	std_logic_vector(15 downto 0) := x"0000"; 
		D		: in 	std_logic_vector(15 downto 0) := x"0000"; 
		O		: out 	std_logic_vector(31 downto 0) ;
		CLK		: in 	std_logic ; 
		CE		: in 	std_logic := 'H' ; 
		IRSTTOP 	: in 	std_logic := 'L' ; 
	    	IRSTBOT 	: in 	std_logic := 'L' ;  
		ORSTTOP 	: in 	std_logic := 'L' ; 
		ORSTBOT 	: in 	std_logic := 'L' ; 
		AHOLD 		: in	std_logic := 'L' ; 
		BHOLD		: in 	std_logic := 'L' ; 
		CHOLD		: in 	std_logic := 'L' ; 
		DHOLD		: in 	std_logic := 'L' ; 
		OHOLDTOP	: in 	std_logic := 'L' ; 
		OHOLDBOT	: in 	std_logic := 'L' ; 
		OLOADTOP	: in	std_logic := 'L' ; 
		OLOADBOT	: in 	std_logic := 'L' ; 
		ADDSUBTOP	: in 	std_logic := 'L' ; 
		ADDSUBBOT	: in 	std_logic := 'L' ;
		CO		: out 	std_logic ;
		CI		: in 	std_logic := 'L' ;  
		ACCUMCI		: in 	std_logic := 'L' ; 
		ACCUMCO        	: out 	std_logic ;
		SIGNEXTIN	: in	std_logic ; 
		SIGNEXTOUT      : out 	std_logic  				
	); 
	attribute VITAL_LEVEL0 of			    
    SB_MAC16  : entity is true;

end SB_MAC16;
	
architecture SB_MAC16_V of SB_MAC16 is
attribute VITAL_LEVEL0 of
SB_MAC16_V : architecture is true; 
	
	signal  Q_zd  : std_logic_vector(31 downto 0)  := (others => 'X');	
	  signal QCO_zd :	 std_ulogic :='X';    
	  signal QACCUMCO_zd :std_ulogic :='X'; 
	  signal SIGNEXTOUT_zd :	 std_ulogic :='X'; 
	signal	A_ipd		: std_logic_vector(15 downto 0)  := (others => 'X');
	signal	B_ipd		:  std_logic_vector(15 downto 0)  := (others => 'X');
	signal	C_ipd		: std_logic_vector(15 downto 0)  := (others => 'X');
	signal	D_ipd		:  std_logic_vector(15 downto 0)  := (others => 'X');
	signal	CLK_ipd		: std_ulogic :='X'; 
	signal	CE_ipd		: std_ulogic :='X';
	signal	IRSTTOP_ipd 	: std_ulogic :='X'; 
	 signal   IRSTBOT_ipd 	: std_ulogic :='X';  
	signal	ORSTTOP_ipd 	: std_ulogic :='X'; 
	signal	ORSTBOT_ipd 	: std_ulogic :='X'; 
	signal	AHOLD_ipd 		:std_ulogic :='X';
	signal	BHOLD_ipd		: std_ulogic :='X'; 
	signal	CHOLD_ipd		: std_ulogic :='X'; 
	signal	DHOLD_ipd		: std_ulogic :='X'; 
	signal	OHOLDTOP_ipd	: std_ulogic :='X'; 
	signal	OHOLDBOT_ipd	: std_ulogic :='X'; 
	signal	OLOADTOP_ipd	:std_ulogic :='X';
	signal	OLOADBOT_ipd	: std_ulogic :='X'; 
	signal	ADDSUBTOP_ipd	: std_ulogic :='X'; 
	signal	ADDSUBBOT_ipd	: std_ulogic :='X';
	signal	CI_ipd		: std_ulogic :='X'; 
	signal	ACCUMCI_ipd		: std_ulogic :='X';
	signal	SIGNEXTIN_ipd	: std_ulogic :='X';	    		  
	-- MULT8/16 which is the check1 so ignore here	


	component mac16_physical is 
	port  (
	 	CLK				: in	std_logic ; 
	 	IHRST				: in	std_logic ;
	 	ILRST				: in	std_logic ;
	 	OHRST				: in	std_logic ;
	 	OLRST				: in	std_logic ;
	 	A 				: in	std_logic_vector (15 downto 0);
	 	B 				: in	std_logic_vector (15 downto 0);
	 	C 				: in	std_logic_vector (15 downto 0);
	 	D 				: in	std_logic_vector (15 downto 0);
	    	CBIT				: in	std_logic_vector (24 downto 0);
	    	AHLD				: in	std_logic ;
	 	BHLD				: in	std_logic ;
	 	CHLD				: in	std_logic ;
	 	DHLD				: in	std_logic ;
	 	OHHLD				: in	std_logic ;
	 	OLHLD				: in	std_logic ;
		OHADS				: in	std_logic ;
	 	OLADS				: in	std_logic ;
	 	OHLDA				: in	std_logic ;
	 	OLLDA				: in	std_logic ;
	 	CICAS				: in	std_logic ;
	 	CI				: in	std_logic ;
	 	SIGNEXTIN			: in	std_logic ;
	 	SIGNEXTOUT			: out	std_logic ;
	 	COCAS				: out	std_logic ;
	 	CO				: out 	std_logic ;
	 	O				: out	std_logic_vector (31 downto 0)	
    	);
	end component; 


	--  for generics 
	signal neg_trig				: std_logic ; 	
	 signal cbitss_inreg			: std_logic_vector(3 downto 0);		    
	signal cbitss_mpyreg			: std_logic_vector(3 downto 0);		   
	signal cbitss_topmac 			: std_logic_vector(6 downto 0);		   
	signal cbitss_botmac 			: std_logic_vector(6 downto 0);		   
	signal cbitss_sign			: std_logic_vector(2 downto 0);		   	
	signal cbitss 				: std_logic_vector (24 downto 0);
	--
	signal  CLK_g , intCLK			: std_logic ; 


begin 

	 	 SIGNEXTOUT	<= SIGNEXTOUT_zd;
	 	-- ACCUMCO		<= ACCUMCO_zd;
	 	-- CO			<= CO_zd;
  WireDelay : block
  begin
    A_DELAY : for i in 15 downto 0 generate
       VitalWireDelay (A_ipd(i), A(i), tipd_A(i));
    end generate A_DELAY;  
    B_DELAY : for i in 15 downto 0 generate
       VitalWireDelay (B_ipd(i), B(i), tipd_B(i));
    end generate B_DELAY;
    C_DELAY : for i in 15 downto 0 generate
       VitalWireDelay (C_ipd(i), C(i), tipd_C(i));
    end generate C_DELAY;
    D_DELAY : for i in 15 downto 0 generate
       VitalWireDelay (D_ipd(i), D(i), tipd_D(i));
    end generate D_DELAY;	
	VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
	VitalWireDelay (CE_ipd, CE_ipd, tipd_CE);
	VitalWireDelay (IRSTTOP_ipd, IRSTTOP, tipd_IRSTTOP);
	VitalWireDelay (IRSTBOT_ipd, IRSTBOT, tipd_IRSTBOT);
	VitalWireDelay (ORSTBOT_ipd, ORSTBOT, tipd_ORSTBOT);
	VitalWireDelay (ORSTTOP_ipd, ORSTTOP, tipd_ORSTTOP);
	VitalWireDelay (AHOLD_ipd, AHOLD, tipd_AHOLD);
	VitalWireDelay (BHOLD_ipd, BHOLD, tipd_BHOLD);
	VitalWireDelay (CHOLD_ipd, CHOLD, tipd_CHOLD);
	VitalWireDelay (DHOLD_ipd, DHOLD, tipd_DHOLD);
	VitalWireDelay (OHOLDTOP_ipd, OHOLDTOP, tipd_OHOLDTOP);
	VitalWireDelay (OHOLDBOT_ipd, OHOLDBOT, tipd_OHOLDBOT);
	VitalWireDelay (OLOADTOP_ipd, OLOADTOP, tipd_OLOADTOP);
	VitalWireDelay (OLOADBOT_ipd, OLOADBOT, tipd_OLOADBOT);
	VitalWireDelay (ADDSUBTOP_ipd, ADDSUBTOP, tipd_ADDSUBTOP);
	VitalWireDelay (ADDSUBBOT_ipd, ADDSUBBOT, tipd_ADDSUBBOT);
	VitalWireDelay (CI_ipd, CI, tipd_CI);
	VitalWireDelay (ACCUMCI_ipd, ACCUMCI, tipd_ACCUMCI);
	VitalWireDelay (SIGNEXTIN_ipd, SIGNEXTIN, tipd_SIGNEXTIN);
end block;


	
	cbitss_inreg 	<= TO_STDLOGICVECTOR( D_REG & B_REG & A_REG & C_REG ); 
    	cbitss_mpyreg   	<= TO_STDLOGICVECTOR( PIPELINE_16x16_MULT_REG2 & PIPELINE_16x16_MULT_REG1 & BOT_8x8_MULT_REG & TOP_8x8_MULT_REG);
    	cbitss_topmac	<= TO_STDLOGICVECTOR( TOPADDSUB_CARRYSELECT & TOPADDSUB_UPPERINPUT & TOPADDSUB_LOWERINPUT & TOPOUTPUT_SELECT );
    	cbitss_botmac	<= TO_STDLOGICVECTOR( BOTADDSUB_CARRYSELECT & BOTADDSUB_UPPERINPUT & BOTADDSUB_LOWERINPUT & BOTOUTPUT_SELECT );
	cbitss_sign	<= TO_STDLOGICVECTOR( B_SIGNED & A_SIGNED & MODE_8x8); 
	cbitss 	  	<= (cbitss_sign & cbitss_botmac & cbitss_topmac & cbitss_mpyreg & cbitss_inreg); 

	---Logic section ---
  	CLK_g <= CLK_ipd and  CE_ipd ;  		   -- CE=0 disables entire clock  
   	intCLK <= (CLK_g xor neg_trig);		   -- Clock Polarity control  
	
	
VITALBehavior : process(	A_ipd,B_ipd,C_ipd,D_ipd,CLK_ipd	,CE_ipd,IRSTTOP_ipd,IRSTBOT_ipd, ORSTTOP_ipd,ORSTBOT_ipd,AHOLD_ipd,BHOLD_ipd,CHOLD_ipd,
DHOLD_ipd,OHOLDTOP_ipd, OHOLDBOT_ipd,OLOADTOP_ipd,OLOADBOT_ipd,ADDSUBTOP_ipd,ADDSUBBOT_ipd,CI_ipd,ACCUMCI_ipd,SIGNEXTIN_ipd,Q_zd,QCO_zd,QACCUMCO_zd,SIGNEXTOUT_zd)

       variable Tviol_A0_CLK_posedge : std_logic := '0';
       variable Tviol_A1_CLK_posedge : std_logic := '0';
       variable Tviol_A2_CLK_posedge : std_logic := '0';
       variable Tviol_A3_CLK_posedge : std_logic := '0';
       variable Tviol_A4_CLK_posedge : std_logic := '0';
       variable Tviol_A5_CLK_posedge : std_logic := '0';
       variable Tviol_A6_CLK_posedge : std_logic := '0';
       variable Tviol_A7_CLK_posedge : std_logic := '0';
	   variable Tviol_A8_CLK_posedge : std_logic := '0';
	   variable Tviol_A9_CLK_posedge : std_logic := '0';
	   variable Tviol_A10_CLK_posedge : std_logic := '0';
	   variable Tviol_A11_CLK_posedge : std_logic := '0';
	   variable Tviol_A12_CLK_posedge : std_logic := '0';
	   variable Tviol_A13_CLK_posedge : std_logic := '0';
	   variable Tviol_A14_CLK_posedge : std_logic := '0';
	   variable Tviol_A15_CLK_posedge : std_logic := '0';

       variable Tmkr_A0_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_A1_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_A2_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_A3_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_A4_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_A5_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_A6_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_A7_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_A8_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_A9_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_A10_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_A11_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_A12_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_A13_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_A14_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_A15_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;	 
	   
	   variable Tviol_B0_CLK_posedge : std_logic := '0';
       variable Tviol_B1_CLK_posedge : std_logic := '0';
       variable Tviol_B2_CLK_posedge : std_logic := '0';
       variable Tviol_B3_CLK_posedge : std_logic := '0';
       variable Tviol_B4_CLK_posedge : std_logic := '0';
       variable Tviol_B5_CLK_posedge : std_logic := '0';
       variable Tviol_B6_CLK_posedge : std_logic := '0';
       variable Tviol_B7_CLK_posedge : std_logic := '0';
	   variable Tviol_B8_CLK_posedge : std_logic := '0';
	   variable Tviol_B9_CLK_posedge : std_logic := '0';
	   variable Tviol_B10_CLK_posedge : std_logic := '0';
	   variable Tviol_B11_CLK_posedge : std_logic := '0';
	   variable Tviol_B12_CLK_posedge : std_logic := '0';
	   variable Tviol_B13_CLK_posedge : std_logic := '0';
	   variable Tviol_B14_CLK_posedge : std_logic := '0';
	   variable Tviol_B15_CLK_posedge : std_logic := '0';

       variable Tmkr_B0_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_B1_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_B2_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_B3_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_B4_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_B5_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_B6_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_B7_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_B8_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_B9_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_B10_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_B11_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_B12_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_B13_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_B14_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_B15_CLK_posedge : VitalTimingDataType := VitalTimingDataInit; 	
	   
	     variable Tviol_C0_CLK_posedge : std_logic := '0';
       variable Tviol_C1_CLK_posedge : std_logic := '0';
       variable Tviol_C2_CLK_posedge : std_logic := '0';
       variable Tviol_C3_CLK_posedge : std_logic := '0';
       variable Tviol_C4_CLK_posedge : std_logic := '0';
       variable Tviol_C5_CLK_posedge : std_logic := '0';
       variable Tviol_C6_CLK_posedge : std_logic := '0';
       variable Tviol_C7_CLK_posedge : std_logic := '0';
	   variable Tviol_C8_CLK_posedge : std_logic := '0';
	   variable Tviol_C9_CLK_posedge : std_logic := '0';
	   variable Tviol_C10_CLK_posedge : std_logic := '0';
	   variable Tviol_C11_CLK_posedge : std_logic := '0';
	   variable Tviol_C12_CLK_posedge : std_logic := '0';
	   variable Tviol_C13_CLK_posedge : std_logic := '0';
	   variable Tviol_C14_CLK_posedge : std_logic := '0';
	   variable Tviol_C15_CLK_posedge : std_logic := '0';

       variable Tmkr_C0_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_C1_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_C2_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_C3_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_C4_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_C5_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_C6_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_C7_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_C8_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_C9_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_C10_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_C11_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_C12_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_C13_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_C14_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_C15_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;	  
	   
	   
	   variable Tviol_D0_CLK_posedge : std_logic := '0';
       variable Tviol_D1_CLK_posedge : std_logic := '0';
       variable Tviol_D2_CLK_posedge : std_logic := '0';
       variable Tviol_D3_CLK_posedge : std_logic := '0';
       variable Tviol_D4_CLK_posedge : std_logic := '0';
       variable Tviol_D5_CLK_posedge : std_logic := '0';
       variable Tviol_D6_CLK_posedge : std_logic := '0';
       variable Tviol_D7_CLK_posedge : std_logic := '0';
	   variable Tviol_D8_CLK_posedge : std_logic := '0';
	   variable Tviol_D9_CLK_posedge : std_logic := '0';
	   variable Tviol_D10_CLK_posedge : std_logic := '0';
	   variable Tviol_D11_CLK_posedge : std_logic := '0';
	   variable Tviol_D12_CLK_posedge : std_logic := '0';
	   variable Tviol_D13_CLK_posedge : std_logic := '0';
	   variable Tviol_D14_CLK_posedge : std_logic := '0';
	   variable Tviol_D15_CLK_posedge : std_logic := '0';

       variable Tmkr_D0_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_D1_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_D2_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_D3_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_D4_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_D5_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_D6_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_D7_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_D8_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_D9_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_D10_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_D11_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_D12_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_D13_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_D14_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   variable Tmkr_D15_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	   
	   variable Tviol_AHOLD_CLK_posedge : std_logic := '0'; 
	   variable Tmkr_AHOLD_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;  
	   variable Tviol_BHOLD_CLK_posedge : std_logic := '0'; 
	   variable Tmkr_BHOLD_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;  
	   
	   variable Tviol_CHOLD_CLK_posedge : std_logic := '0'; 
	   variable Tmkr_CHOLD_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;  
	   
	   variable Tviol_DHOLD_CLK_posedge : std_logic := '0'; 
	   variable Tmkr_DHOLD_CLK_posedge : VitalTimingDataType := VitalTimingDataInit; 	
	   
	    variable Tviol_ADDSUBTOP_CLK_posedge : std_logic := '0'; 
	   variable Tmkr_ADDSUBTOP_CLK_posedge : VitalTimingDataType := VitalTimingDataInit; 
	   
	    variable Tviol_ADDSUBBOT_CLK_posedge : std_logic := '0'; 
	   variable Tmkr_ADDSUBBOT_CLK_posedge : VitalTimingDataType := VitalTimingDataInit; 
	   
	    variable Tviol_OHOLDTOP_CLK_posedge : std_logic := '0'; 
	   variable Tmkr_OHOLDTOP_CLK_posedge : VitalTimingDataType := VitalTimingDataInit; 
	   
	   	   variable Tviol_OHOLDBOT_CLK_posedge : std_logic := '0'; 
	   variable Tmkr_OHOLDBOT_CLK_posedge : VitalTimingDataType := VitalTimingDataInit; 
	   
	   	   variable Tviol_OLOADTOP_CLK_posedge : std_logic := '0'; 
	   variable Tmkr_OLOADTOP_CLK_posedge : VitalTimingDataType := VitalTimingDataInit; 
	   
	   	   variable Tviol_OLOADBOT_CLK_posedge : std_logic := '0'; 
	   variable Tmkr_OLOADBOT_CLK_posedge : VitalTimingDataType := VitalTimingDataInit; 

	   	   	variable Tviol_CI_CLK_posedge : std_logic := '0'; 
	   variable Tmkr_CI_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;  
	   
	   variable Tviol_ACCUMCI_CLK_posedge : std_logic := '0'; 
	   variable Tmkr_ACCUMCI_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;  
	   
	           variable PViol_CLK : std_logic := '0';

        variable PInfo_CLK : VitalPeriodDataType := VitalPeriodDataInit;	
		
		variable Tviol_IRSTTOP_CLK_posedge: std_logic := '0';
		variable Tmkr_IRSTTOP_CLK_posedge : VitalTimingDataType := VitalTimingDataInit; 
		variable Tviol_IRSTBOT_CLK_posedge: std_logic := '0';
		variable Tmkr_IRSTBOT_CLK_posedge : VitalTimingDataType := VitalTimingDataInit; 
		variable Tviol_ORSTTOP_CLK_posedge: std_logic := '0';
		variable Tmkr_ORSTTOP_CLK_posedge : VitalTimingDataType := VitalTimingDataInit; 
		variable Tviol_ORSTBOT_CLK_posedge: std_logic := '0';
		variable Tmkr_ORSTBOT_CLK_posedge : VitalTimingDataType := VitalTimingDataInit; 	
		
		variable Tviol_IRSTTOP_CLK_negedge: std_logic := '0';
		variable Tmkr_IRSTTOP_CLK_negedge : VitalTimingDataType := VitalTimingDataInit; 
		variable Tviol_IRSTBOT_CLK_negedge: std_logic := '0';
		variable Tmkr_IRSTBOT_CLK_negedge : VitalTimingDataType := VitalTimingDataInit; 
		variable Tviol_ORSTTOP_CLK_negedge: std_logic := '0';
		variable Tmkr_ORSTTOP_CLK_negedge : VitalTimingDataType := VitalTimingDataInit; 
		variable Tviol_ORSTBOT_CLK_negedge: std_logic := '0';
		variable Tmkr_ORSTBOT_CLK_negedge : VitalTimingDataType := VitalTimingDataInit;
		
		--variable O_GlitchData  : VitalGlitchDataArrayType (31 downto 0);
		
		
begin 

    if (TimingChecksOn) then
      VitalSetupHoldCheck (
        Violation      => Tviol_A0_CLK_posedge,
        TimingData     => Tmkr_A0_CLK_posedge,
        TestSignal     => A_ipd(0),
        TestSignalName => "A(0)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_A_CLK_posedge_posedge(0),
        SetupLow       => tsetup_A_CLK_negedge_posedge(0),
        HoldLow        => thold_A_CLK_posedge_posedge(0),
        HoldHigh       => thold_A_CLK_negedge_posedge(0),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	 
		    VitalSetupHoldCheck (
        Violation      => Tviol_A1_CLK_posedge,
        TimingData     => Tmkr_A1_CLK_posedge,
        TestSignal     => A_ipd(1),
        TestSignalName => "A(1)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_A_CLK_posedge_posedge(1),
        SetupLow       => tsetup_A_CLK_negedge_posedge(1),
        HoldLow        => thold_A_CLK_posedge_posedge(1),
        HoldHigh       => thold_A_CLK_negedge_posedge(1),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_A2_CLK_posedge,
        TimingData     => Tmkr_A2_CLK_posedge,
        TestSignal     => A_ipd(2),
        TestSignalName => "A(2)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_A_CLK_posedge_posedge(2),
        SetupLow       => tsetup_A_CLK_negedge_posedge(2),
        HoldLow        => thold_A_CLK_posedge_posedge(2),
        HoldHigh       => thold_A_CLK_negedge_posedge(2),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_A3_CLK_posedge,
        TimingData     => Tmkr_A3_CLK_posedge,
        TestSignal     => A_ipd(3),
        TestSignalName => "A(3)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_A_CLK_posedge_posedge(3),
        SetupLow       => tsetup_A_CLK_negedge_posedge(3),
        HoldLow        => thold_A_CLK_posedge_posedge(3),
        HoldHigh       => thold_A_CLK_negedge_posedge(3),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_A4_CLK_posedge,
        TimingData     => Tmkr_A4_CLK_posedge,
        TestSignal     => A_ipd(4),
        TestSignalName => "A(4)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_A_CLK_posedge_posedge(4),
        SetupLow       => tsetup_A_CLK_negedge_posedge(4),
        HoldLow        => thold_A_CLK_posedge_posedge(4),
        HoldHigh       => thold_A_CLK_negedge_posedge(4),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_A5_CLK_posedge,
        TimingData     => Tmkr_A5_CLK_posedge,
        TestSignal     => A_ipd(5),
        TestSignalName => "A(5)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_A_CLK_posedge_posedge(5),
        SetupLow       => tsetup_A_CLK_negedge_posedge(5),
        HoldLow        => thold_A_CLK_posedge_posedge(5),
        HoldHigh       => thold_A_CLK_negedge_posedge(5),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_A6_CLK_posedge,
        TimingData     => Tmkr_A6_CLK_posedge,
        TestSignal     => A_ipd(6),
        TestSignalName => "A(6)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_A_CLK_posedge_posedge(6),
        SetupLow       => tsetup_A_CLK_negedge_posedge(6),
        HoldLow        => thold_A_CLK_posedge_posedge(6),
        HoldHigh       => thold_A_CLK_negedge_posedge(6),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_A7_CLK_posedge,
        TimingData     => Tmkr_A7_CLK_posedge,
        TestSignal     => A_ipd(7),
        TestSignalName => "A(7)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_A_CLK_posedge_posedge(7),
        SetupLow       => tsetup_A_CLK_negedge_posedge(7),
        HoldLow        => thold_A_CLK_posedge_posedge(7),
        HoldHigh       => thold_A_CLK_negedge_posedge(7),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_A8_CLK_posedge,
        TimingData     => Tmkr_A8_CLK_posedge,
        TestSignal     => A_ipd(8),
        TestSignalName => "A(8)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_A_CLK_posedge_posedge(8),
        SetupLow       => tsetup_A_CLK_negedge_posedge(8),
        HoldLow        => thold_A_CLK_posedge_posedge(8),
        HoldHigh       => thold_A_CLK_negedge_posedge(8),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_A9_CLK_posedge,
        TimingData     => Tmkr_A9_CLK_posedge,
        TestSignal     => A_ipd(9),
        TestSignalName => "A(9)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_A_CLK_posedge_posedge(9),
        SetupLow       => tsetup_A_CLK_negedge_posedge(9),
        HoldLow        => thold_A_CLK_posedge_posedge(9),
        HoldHigh       => thold_A_CLK_negedge_posedge(9),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_A10_CLK_posedge,
        TimingData     => Tmkr_A10_CLK_posedge,
        TestSignal     => A_ipd(10),
        TestSignalName => "A(10)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_A_CLK_posedge_posedge(10),
        SetupLow       => tsetup_A_CLK_negedge_posedge(10),
        HoldLow        => thold_A_CLK_posedge_posedge(10),
        HoldHigh       => thold_A_CLK_negedge_posedge(10),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_A11_CLK_posedge,
        TimingData     => Tmkr_A11_CLK_posedge,
        TestSignal     => A_ipd(11),
        TestSignalName => "A(11)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_A_CLK_posedge_posedge(11),
        SetupLow       => tsetup_A_CLK_negedge_posedge(11),
        HoldLow        => thold_A_CLK_posedge_posedge(11),
        HoldHigh       => thold_A_CLK_negedge_posedge(11),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_A12_CLK_posedge,
        TimingData     => Tmkr_A12_CLK_posedge,
        TestSignal     => A_ipd(12),
        TestSignalName => "A(12)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_A_CLK_posedge_posedge(12),
        SetupLow       => tsetup_A_CLK_negedge_posedge(12),
        HoldLow        => thold_A_CLK_posedge_posedge(12),
        HoldHigh       => thold_A_CLK_negedge_posedge(12),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_A13_CLK_posedge,
        TimingData     => Tmkr_A13_CLK_posedge,
        TestSignal     => A_ipd(13),
        TestSignalName => "A(13)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_A_CLK_posedge_posedge(13),
        SetupLow       => tsetup_A_CLK_negedge_posedge(13),
        HoldLow        => thold_A_CLK_posedge_posedge(13),
        HoldHigh       => thold_A_CLK_negedge_posedge(13),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_A14_CLK_posedge,
        TimingData     => Tmkr_A14_CLK_posedge,
        TestSignal     => A_ipd(14),
        TestSignalName => "A(14)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_A_CLK_posedge_posedge(14),
        SetupLow       => tsetup_A_CLK_negedge_posedge(14),
        HoldLow        => thold_A_CLK_posedge_posedge(14),
        HoldHigh       => thold_A_CLK_negedge_posedge(14),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_A15_CLK_posedge,
        TimingData     => Tmkr_A15_CLK_posedge,
        TestSignal     => A_ipd(15),
        TestSignalName => "A(15)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_A_CLK_posedge_posedge(15),
        SetupLow       => tsetup_A_CLK_negedge_posedge(15),
        HoldLow        => thold_A_CLK_posedge_posedge(15),
        HoldHigh       => thold_A_CLK_negedge_posedge(15),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		 
		    
		VitalSetupHoldCheck (
        Violation      => Tviol_B0_CLK_posedge,
        TimingData     => Tmkr_B0_CLK_posedge,
        TestSignal     => B_ipd(0),
        TestSignalName => "B(0)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_B_CLK_posedge_posedge(0),
        SetupLow       => tsetup_B_CLK_negedge_posedge(0),
        HoldLow        => thold_B_CLK_posedge_posedge(0),
        HoldHigh       => thold_B_CLK_negedge_posedge(0),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	 
		   VitalSetupHoldCheck (
        Violation      => Tviol_B1_CLK_posedge,
        TimingData     => Tmkr_B1_CLK_posedge,
        TestSignal     => B_ipd(1),
        TestSignalName => "B(1)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_B_CLK_posedge_posedge(1),
        SetupLow       => tsetup_B_CLK_negedge_posedge(1),
        HoldLow        => thold_B_CLK_posedge_posedge(1),
        HoldHigh       => thold_B_CLK_negedge_posedge(1),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_B2_CLK_posedge,
        TimingData     => Tmkr_B2_CLK_posedge,
        TestSignal     => B_ipd(2),
        TestSignalName => "B(2)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_B_CLK_posedge_posedge(2),
        SetupLow       => tsetup_B_CLK_negedge_posedge(2),
        HoldLow        => thold_B_CLK_posedge_posedge(2),
        HoldHigh       => thold_B_CLK_negedge_posedge(2),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_B3_CLK_posedge,
        TimingData     => Tmkr_B3_CLK_posedge,
        TestSignal     => B_ipd(3),
        TestSignalName => "B(3)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_B_CLK_posedge_posedge(3),
        SetupLow       => tsetup_B_CLK_negedge_posedge(3),
        HoldLow        => thold_B_CLK_posedge_posedge(3),
        HoldHigh       => thold_B_CLK_negedge_posedge(3),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_B4_CLK_posedge,
        TimingData     => Tmkr_B4_CLK_posedge,
        TestSignal     => B_ipd(4),
        TestSignalName => "B(4)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_B_CLK_posedge_posedge(4),
        SetupLow       => tsetup_B_CLK_negedge_posedge(4),
        HoldLow        => thold_B_CLK_posedge_posedge(4),
        HoldHigh       => thold_B_CLK_negedge_posedge(4),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_B5_CLK_posedge,
        TimingData     => Tmkr_B5_CLK_posedge,
        TestSignal     => B_ipd(5),
        TestSignalName => "B(5)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_B_CLK_posedge_posedge(5),
        SetupLow       => tsetup_B_CLK_negedge_posedge(5),
        HoldLow        => thold_B_CLK_posedge_posedge(5),
        HoldHigh       => thold_B_CLK_negedge_posedge(5),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_B6_CLK_posedge,
        TimingData     => Tmkr_B6_CLK_posedge,
        TestSignal     => B_ipd(6),
        TestSignalName => "B(6)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_B_CLK_posedge_posedge(6),
        SetupLow       => tsetup_B_CLK_negedge_posedge(6),
        HoldLow        => thold_B_CLK_posedge_posedge(6),
        HoldHigh       => thold_B_CLK_negedge_posedge(6),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_B7_CLK_posedge,
        TimingData     => Tmkr_B7_CLK_posedge,
        TestSignal     => B_ipd(7),
        TestSignalName => "B(7)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_B_CLK_posedge_posedge(7),
        SetupLow       => tsetup_B_CLK_negedge_posedge(7),
        HoldLow        => thold_B_CLK_posedge_posedge(7),
        HoldHigh       => thold_B_CLK_negedge_posedge(7),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_B8_CLK_posedge,
        TimingData     => Tmkr_B8_CLK_posedge,
        TestSignal     => B_ipd(8),
        TestSignalName => "B(8)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_B_CLK_posedge_posedge(8),
        SetupLow       => tsetup_B_CLK_negedge_posedge(8),
        HoldLow        => thold_B_CLK_posedge_posedge(8),
        HoldHigh       => thold_B_CLK_negedge_posedge(8),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_B9_CLK_posedge,
        TimingData     => Tmkr_B9_CLK_posedge,
        TestSignal     => B_ipd(9),
        TestSignalName => "B(9)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_B_CLK_posedge_posedge(9),
        SetupLow       => tsetup_B_CLK_negedge_posedge(9),
        HoldLow        => thold_B_CLK_posedge_posedge(9),
        HoldHigh       => thold_B_CLK_negedge_posedge(9),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_B10_CLK_posedge,
        TimingData     => Tmkr_B10_CLK_posedge,
        TestSignal     => B_ipd(10),
        TestSignalName => "B(10)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_B_CLK_posedge_posedge(10),
        SetupLow       => tsetup_B_CLK_negedge_posedge(10),
        HoldLow        => thold_B_CLK_posedge_posedge(10),
        HoldHigh       => thold_B_CLK_negedge_posedge(10),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_B11_CLK_posedge,
        TimingData     => Tmkr_B11_CLK_posedge,
        TestSignal     => B_ipd(11),
        TestSignalName => "B(11)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_B_CLK_posedge_posedge(11),
        SetupLow       => tsetup_B_CLK_negedge_posedge(11),
        HoldLow        => thold_B_CLK_posedge_posedge(11),
        HoldHigh       => thold_B_CLK_negedge_posedge(11),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_B12_CLK_posedge,
        TimingData     => Tmkr_B12_CLK_posedge,
        TestSignal     => B_ipd(12),
        TestSignalName => "B(12)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_B_CLK_posedge_posedge(12),
        SetupLow       => tsetup_B_CLK_negedge_posedge(12),
        HoldLow        => thold_B_CLK_posedge_posedge(12),
        HoldHigh       => thold_B_CLK_negedge_posedge(12),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_B13_CLK_posedge,
        TimingData     => Tmkr_B13_CLK_posedge,
        TestSignal     => B_ipd(13),
        TestSignalName => "B(13)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_B_CLK_posedge_posedge(13),
        SetupLow       => tsetup_B_CLK_negedge_posedge(13),
        HoldLow        => thold_B_CLK_posedge_posedge(13),
        HoldHigh       => thold_B_CLK_negedge_posedge(13),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_B14_CLK_posedge,
        TimingData     => Tmkr_B14_CLK_posedge,
        TestSignal     => B_ipd(14),
        TestSignalName => "B(14)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_B_CLK_posedge_posedge(14),
        SetupLow       => tsetup_B_CLK_negedge_posedge(14),
        HoldLow        => thold_B_CLK_posedge_posedge(14),
        HoldHigh       => thold_B_CLK_negedge_posedge(14),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_B15_CLK_posedge,
        TimingData     => Tmkr_B15_CLK_posedge,
        TestSignal     => B_ipd(15),
        TestSignalName => "B(15)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_B_CLK_posedge_posedge(15),
        SetupLow       => tsetup_B_CLK_negedge_posedge(15),
        HoldLow        => thold_B_CLK_posedge_posedge(15),
        HoldHigh       => thold_B_CLK_negedge_posedge(15),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	 
		
		
		    VitalSetupHoldCheck (
        Violation      => Tviol_AHOLD_CLK_posedge,
        TimingData     => Tmkr_AHOLD_CLK_posedge,
        TestSignal     => AHOLD_ipd,
        TestSignalName => "AHOLD",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_AHOLD_CLK_posedge_posedge,
        SetupLow       => tsetup_AHOLD_CLK_negedge_posedge,
        HoldLow        => thold_AHOLD_CLK_posedge_posedge,
        HoldHigh       => thold_AHOLD_CLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	  
		
		
		    VitalSetupHoldCheck (
        Violation      => Tviol_BHOLD_CLK_posedge,
        TimingData     => Tmkr_BHOLD_CLK_posedge,
        TestSignal     => BHOLD_ipd,
        TestSignalName => "BHOLD",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_BHOLD_CLK_posedge_posedge,
        SetupLow       => tsetup_BHOLD_CLK_negedge_posedge,
        HoldLow        => thold_BHOLD_CLK_posedge_posedge,
        HoldHigh       => thold_BHOLD_CLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		
		
		
		VitalSetupHoldCheck (
        Violation      => Tviol_C0_CLK_posedge,
        TimingData     => Tmkr_C0_CLK_posedge,
        TestSignal     => C_ipd(0),
        TestSignalName => "C(0)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_C_CLK_posedge_posedge(0),
        SetupLow       => tsetup_C_CLK_negedge_posedge(0),
        HoldLow        => thold_C_CLK_posedge_posedge(0),
        HoldHigh       => thold_C_CLK_negedge_posedge(0),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	 
		    VitalSetupHoldCheck (
        Violation      => Tviol_C1_CLK_posedge,
        TimingData     => Tmkr_C1_CLK_posedge,
        TestSignal     => C_ipd(1),
        TestSignalName => "C(1)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_C_CLK_posedge_posedge(1),
        SetupLow       => tsetup_C_CLK_negedge_posedge(1),
        HoldLow        => thold_C_CLK_posedge_posedge(1),
        HoldHigh       => thold_C_CLK_negedge_posedge(1),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_C2_CLK_posedge,
        TimingData     => Tmkr_C2_CLK_posedge,
        TestSignal     => C_ipd(2),
        TestSignalName => "C(2)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_C_CLK_posedge_posedge(2),
        SetupLow       => tsetup_C_CLK_negedge_posedge(2),
        HoldLow        => thold_C_CLK_posedge_posedge(2),
        HoldHigh       => thold_C_CLK_negedge_posedge(2),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_C3_CLK_posedge,
        TimingData     => Tmkr_C3_CLK_posedge,
        TestSignal     => C_ipd(3),
        TestSignalName => "C(3)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_C_CLK_posedge_posedge(3),
        SetupLow       => tsetup_C_CLK_negedge_posedge(3),
        HoldLow        => thold_C_CLK_posedge_posedge(3),
        HoldHigh       => thold_C_CLK_negedge_posedge(3),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_C4_CLK_posedge,
        TimingData     => Tmkr_C4_CLK_posedge,
        TestSignal     => C_ipd(4),
        TestSignalName => "C(4)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_C_CLK_posedge_posedge(4),
        SetupLow       => tsetup_C_CLK_negedge_posedge(4),
        HoldLow        => thold_C_CLK_posedge_posedge(4),
        HoldHigh       => thold_C_CLK_negedge_posedge(4),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_C5_CLK_posedge,
        TimingData     => Tmkr_C5_CLK_posedge,
        TestSignal     => C_ipd(5),
        TestSignalName => "C(5)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_C_CLK_posedge_posedge(5),
        SetupLow       => tsetup_C_CLK_negedge_posedge(5),
        HoldLow        => thold_C_CLK_posedge_posedge(5),
        HoldHigh       => thold_C_CLK_negedge_posedge(5),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_C6_CLK_posedge,
        TimingData     => Tmkr_C6_CLK_posedge,
        TestSignal     => C_ipd(6),
        TestSignalName => "C(6)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_C_CLK_posedge_posedge(6),
        SetupLow       => tsetup_C_CLK_negedge_posedge(6),
        HoldLow        => thold_C_CLK_posedge_posedge(6),
        HoldHigh       => thold_C_CLK_negedge_posedge(6),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_C7_CLK_posedge,
        TimingData     => Tmkr_C7_CLK_posedge,
        TestSignal     => C_ipd(7),
        TestSignalName => "C(7)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_C_CLK_posedge_posedge(7),
        SetupLow       => tsetup_C_CLK_negedge_posedge(7),
        HoldLow        => thold_C_CLK_posedge_posedge(7),
        HoldHigh       => thold_C_CLK_negedge_posedge(7),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_C8_CLK_posedge,
        TimingData     => Tmkr_C8_CLK_posedge,
        TestSignal     => C_ipd(8),
        TestSignalName => "C(8)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_C_CLK_posedge_posedge(8),
        SetupLow       => tsetup_C_CLK_negedge_posedge(8),
        HoldLow        => thold_C_CLK_posedge_posedge(8),
        HoldHigh       => thold_C_CLK_negedge_posedge(8),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_C9_CLK_posedge,
        TimingData     => Tmkr_C9_CLK_posedge,
        TestSignal     => C_ipd(9),
        TestSignalName => "C(9)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_C_CLK_posedge_posedge(9),
        SetupLow       => tsetup_C_CLK_negedge_posedge(9),
        HoldLow        => thold_C_CLK_posedge_posedge(9),
        HoldHigh       => thold_C_CLK_negedge_posedge(9),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_C10_CLK_posedge,
        TimingData     => Tmkr_C10_CLK_posedge,
        TestSignal     => C_ipd(10),
        TestSignalName => "C(10)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_C_CLK_posedge_posedge(10),
        SetupLow       => tsetup_C_CLK_negedge_posedge(10),
        HoldLow        => thold_C_CLK_posedge_posedge(10),
        HoldHigh       => thold_C_CLK_negedge_posedge(10),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_C11_CLK_posedge,
        TimingData     => Tmkr_C11_CLK_posedge,
        TestSignal     => C_ipd(11),
        TestSignalName => "C(11)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_C_CLK_posedge_posedge(11),
        SetupLow       => tsetup_C_CLK_negedge_posedge(11),
        HoldLow        => thold_C_CLK_posedge_posedge(11),
        HoldHigh       => thold_C_CLK_negedge_posedge(11),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_C12_CLK_posedge,
        TimingData     => Tmkr_C12_CLK_posedge,
        TestSignal     => C_ipd(12),
        TestSignalName => "C(12)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_C_CLK_posedge_posedge(12),
        SetupLow       => tsetup_C_CLK_negedge_posedge(12),
        HoldLow        => thold_C_CLK_posedge_posedge(12),
        HoldHigh       => thold_C_CLK_negedge_posedge(12),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_C13_CLK_posedge,
        TimingData     => Tmkr_C13_CLK_posedge,
        TestSignal     => C_ipd(13),
        TestSignalName => "C(13)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_C_CLK_posedge_posedge(13),
        SetupLow       => tsetup_C_CLK_negedge_posedge(13),
        HoldLow        => thold_C_CLK_posedge_posedge(13),
        HoldHigh       => thold_C_CLK_negedge_posedge(13),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_C14_CLK_posedge,
        TimingData     => Tmkr_C14_CLK_posedge,
        TestSignal     => C_ipd(14),
        TestSignalName => "C(14)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_C_CLK_posedge_posedge(14),
        SetupLow       => tsetup_C_CLK_negedge_posedge(14),
        HoldLow        => thold_C_CLK_posedge_posedge(14),
        HoldHigh       => thold_C_CLK_negedge_posedge(14),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_C15_CLK_posedge,
        TimingData     => Tmkr_C15_CLK_posedge,
        TestSignal     => C_ipd(15),
        TestSignalName => "C(15)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_C_CLK_posedge_posedge(15),
        SetupLow       => tsetup_C_CLK_negedge_posedge(15),
        HoldLow        => thold_C_CLK_posedge_posedge(15),
        HoldHigh       => thold_C_CLK_negedge_posedge(15),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		 
		
			    
		VitalSetupHoldCheck (
        Violation      => Tviol_D0_CLK_posedge,
        TimingData     => Tmkr_D0_CLK_posedge,
        TestSignal     => D_ipd(0),
        TestSignalName => "D(0)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_D_CLK_posedge_posedge(0),
        SetupLow       => tsetup_D_CLK_negedge_posedge(0),
        HoldLow        => thold_D_CLK_posedge_posedge(0),
        HoldHigh       => thold_D_CLK_negedge_posedge(0),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SD_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	 
		   VitalSetupHoldCheck (
        Violation      => Tviol_D1_CLK_posedge,
        TimingData     => Tmkr_D1_CLK_posedge,
        TestSignal     => D_ipd(1),
        TestSignalName => "D(1)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_D_CLK_posedge_posedge(1),
        SetupLow       => tsetup_D_CLK_negedge_posedge(1),
        HoldLow        => thold_D_CLK_posedge_posedge(1),
        HoldHigh       => thold_D_CLK_negedge_posedge(1),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SD_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_D2_CLK_posedge,
        TimingData     => Tmkr_D2_CLK_posedge,
        TestSignal     => D_ipd(2),
        TestSignalName => "D(2)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_D_CLK_posedge_posedge(2),
        SetupLow       => tsetup_D_CLK_negedge_posedge(2),
        HoldLow        => thold_D_CLK_posedge_posedge(2),
        HoldHigh       => thold_D_CLK_negedge_posedge(2),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SD_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_D3_CLK_posedge,
        TimingData     => Tmkr_D3_CLK_posedge,
        TestSignal     => D_ipd(3),
        TestSignalName => "D(3)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_D_CLK_posedge_posedge(3),
        SetupLow       => tsetup_D_CLK_negedge_posedge(3),
        HoldLow        => thold_D_CLK_posedge_posedge(3),
        HoldHigh       => thold_D_CLK_negedge_posedge(3),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SD_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_D4_CLK_posedge,
        TimingData     => Tmkr_D4_CLK_posedge,
        TestSignal     => D_ipd(4),
        TestSignalName => "D(4)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_D_CLK_posedge_posedge(4),
        SetupLow       => tsetup_D_CLK_negedge_posedge(4),
        HoldLow        => thold_D_CLK_posedge_posedge(4),
        HoldHigh       => thold_D_CLK_negedge_posedge(4),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SD_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_D5_CLK_posedge,
        TimingData     => Tmkr_D5_CLK_posedge,
        TestSignal     => D_ipd(5),
        TestSignalName => "D(5)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_D_CLK_posedge_posedge(5),
        SetupLow       => tsetup_D_CLK_negedge_posedge(5),
        HoldLow        => thold_D_CLK_posedge_posedge(5),
        HoldHigh       => thold_D_CLK_negedge_posedge(5),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SD_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_D6_CLK_posedge,
        TimingData     => Tmkr_D6_CLK_posedge,
        TestSignal     => D_ipd(6),
        TestSignalName => "D(6)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_D_CLK_posedge_posedge(6),
        SetupLow       => tsetup_D_CLK_negedge_posedge(6),
        HoldLow        => thold_D_CLK_posedge_posedge(6),
        HoldHigh       => thold_D_CLK_negedge_posedge(6),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SD_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_D7_CLK_posedge,
        TimingData     => Tmkr_D7_CLK_posedge,
        TestSignal     => D_ipd(7),
        TestSignalName => "D(7)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_D_CLK_posedge_posedge(7),
        SetupLow       => tsetup_D_CLK_negedge_posedge(7),
        HoldLow        => thold_D_CLK_posedge_posedge(7),
        HoldHigh       => thold_D_CLK_negedge_posedge(7),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SD_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_D8_CLK_posedge,
        TimingData     => Tmkr_D8_CLK_posedge,
        TestSignal     => D_ipd(8),
        TestSignalName => "D(8)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_D_CLK_posedge_posedge(8),
        SetupLow       => tsetup_D_CLK_negedge_posedge(8),
        HoldLow        => thold_D_CLK_posedge_posedge(8),
        HoldHigh       => thold_D_CLK_negedge_posedge(8),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SD_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_D9_CLK_posedge,
        TimingData     => Tmkr_D9_CLK_posedge,
        TestSignal     => D_ipd(9),
        TestSignalName => "D(9)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_D_CLK_posedge_posedge(9),
        SetupLow       => tsetup_D_CLK_negedge_posedge(9),
        HoldLow        => thold_D_CLK_posedge_posedge(9),
        HoldHigh       => thold_D_CLK_negedge_posedge(9),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SD_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_D10_CLK_posedge,
        TimingData     => Tmkr_D10_CLK_posedge,
        TestSignal     => D_ipd(10),
        TestSignalName => "D(10)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_D_CLK_posedge_posedge(10),
        SetupLow       => tsetup_D_CLK_negedge_posedge(10),
        HoldLow        => thold_D_CLK_posedge_posedge(10),
        HoldHigh       => thold_D_CLK_negedge_posedge(10),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SD_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_D11_CLK_posedge,
        TimingData     => Tmkr_D11_CLK_posedge,
        TestSignal     => D_ipd(11),
        TestSignalName => "D(11)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_D_CLK_posedge_posedge(11),
        SetupLow       => tsetup_D_CLK_negedge_posedge(11),
        HoldLow        => thold_D_CLK_posedge_posedge(11),
        HoldHigh       => thold_D_CLK_negedge_posedge(11),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SD_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_D12_CLK_posedge,
        TimingData     => Tmkr_D12_CLK_posedge,
        TestSignal     => D_ipd(12),
        TestSignalName => "D(12)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_D_CLK_posedge_posedge(12),
        SetupLow       => tsetup_D_CLK_negedge_posedge(12),
        HoldLow        => thold_D_CLK_posedge_posedge(12),
        HoldHigh       => thold_D_CLK_negedge_posedge(12),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SD_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_D13_CLK_posedge,
        TimingData     => Tmkr_D13_CLK_posedge,
        TestSignal     => D_ipd(13),
        TestSignalName => "D(13)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_D_CLK_posedge_posedge(13),
        SetupLow       => tsetup_D_CLK_negedge_posedge(13),
        HoldLow        => thold_D_CLK_posedge_posedge(13),
        HoldHigh       => thold_D_CLK_negedge_posedge(13),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SD_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_D14_CLK_posedge,
        TimingData     => Tmkr_D14_CLK_posedge,
        TestSignal     => D_ipd(14),
        TestSignalName => "D(14)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_D_CLK_posedge_posedge(14),
        SetupLow       => tsetup_D_CLK_negedge_posedge(14),
        HoldLow        => thold_D_CLK_posedge_posedge(14),
        HoldHigh       => thold_D_CLK_negedge_posedge(14),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SD_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		    VitalSetupHoldCheck (
        Violation      => Tviol_D15_CLK_posedge,
        TimingData     => Tmkr_D15_CLK_posedge,
        TestSignal     => D_ipd(15),
        TestSignalName => "D(15)",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_D_CLK_posedge_posedge(15),
        SetupLow       => tsetup_D_CLK_negedge_posedge(15),
        HoldLow        => thold_D_CLK_posedge_posedge(15),
        HoldHigh       => thold_D_CLK_negedge_posedge(15),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SD_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	   
		
		
		 VitalSetupHoldCheck (
        Violation      => Tviol_CHOLD_CLK_posedge,
        TimingData     => Tmkr_CHOLD_CLK_posedge,
        TestSignal     => CHOLD_ipd,
        TestSignalName => "CHOLD",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_CHOLD_CLK_posedge_posedge,
        SetupLow       => tsetup_CHOLD_CLK_negedge_posedge,
        HoldLow        => thold_CHOLD_CLK_posedge_posedge,
        HoldHigh       => thold_CHOLD_CLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	  
		
		 VitalSetupHoldCheck (
        Violation      => Tviol_DHOLD_CLK_posedge,
        TimingData     => Tmkr_DHOLD_CLK_posedge,
        TestSignal     => DHOLD_ipd,
        TestSignalName => "DHOLD",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_DHOLD_CLK_posedge_posedge,
        SetupLow       => tsetup_DHOLD_CLK_negedge_posedge,
        HoldLow        => thold_DHOLD_CLK_posedge_posedge,
        HoldHigh       => thold_DHOLD_CLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		
		
		 VitalSetupHoldCheck (
        Violation      => Tviol_ADDSUBTOP_CLK_posedge,
        TimingData     => Tmkr_ADDSUBTOP_CLK_posedge,
        TestSignal     => ADDSUBTOP_ipd,
        TestSignalName => "ADDSUBTOP",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_ADDSUBTOP_CLK_posedge_posedge,
        SetupLow       => tsetup_ADDSUBTOP_CLK_negedge_posedge,
        HoldLow        => thold_ADDSUBTOP_CLK_posedge_posedge,
        HoldHigh       => thold_ADDSUBTOP_CLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		
		 VitalSetupHoldCheck (
        Violation      => Tviol_ADDSUBBOT_CLK_posedge,
        TimingData     => Tmkr_ADDSUBBOT_CLK_posedge,
        TestSignal     => ADDSUBBOT_ipd,
        TestSignalName => "ADDSUBBOT",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_ADDSUBBOT_CLK_posedge_posedge,
        SetupLow       => tsetup_ADDSUBBOT_CLK_negedge_posedge,
        HoldLow        => thold_ADDSUBBOT_CLK_posedge_posedge,
        HoldHigh       => thold_ADDSUBBOT_CLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		
		 VitalSetupHoldCheck (
        Violation      => Tviol_OHOLDTOP_CLK_posedge,
        TimingData     => Tmkr_OHOLDTOP_CLK_posedge,
        TestSignal     => OHOLDTOP_ipd,
        TestSignalName => "OHOLDTOP",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_OHOLDTOP_CLK_posedge_posedge,
        SetupLow       => tsetup_OHOLDTOP_CLK_negedge_posedge,
        HoldLow        => thold_OHOLDTOP_CLK_posedge_posedge,
        HoldHigh       => thold_OHOLDTOP_CLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		
		 VitalSetupHoldCheck (
        Violation      => Tviol_OHOLDBOT_CLK_posedge,
        TimingData     => Tmkr_OHOLDBOT_CLK_posedge,
        TestSignal     => OHOLDBOT_ipd,
        TestSignalName => "OHOLDBOT",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_OHOLDBOT_CLK_posedge_posedge,
        SetupLow       => tsetup_OHOLDBOT_CLK_negedge_posedge,
        HoldLow        => thold_OHOLDBOT_CLK_posedge_posedge,
        HoldHigh       => thold_OHOLDBOT_CLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		
		 VitalSetupHoldCheck (
        Violation      => Tviol_OLOADTOP_CLK_posedge,
        TimingData     => Tmkr_OLOADTOP_CLK_posedge,
        TestSignal     => OLOADTOP_ipd,
        TestSignalName => "OLOADTOP",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_OLOADTOP_CLK_posedge_posedge,
        SetupLow       => tsetup_OLOADTOP_CLK_negedge_posedge,
        HoldLow        => thold_OLOADTOP_CLK_posedge_posedge,
        HoldHigh       => thold_OLOADTOP_CLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		
		 VitalSetupHoldCheck (
        Violation      => Tviol_OLOADBOT_CLK_posedge,
        TimingData     => Tmkr_OLOADBOT_CLK_posedge,
        TestSignal     => OLOADBOT_ipd,
        TestSignalName => "OLOADBOT",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_OLOADBOT_CLK_posedge_posedge,
        SetupLow       => tsetup_OLOADBOT_CLK_negedge_posedge,
        HoldLow        => thold_OLOADBOT_CLK_posedge_posedge,
        HoldHigh       => thold_OLOADBOT_CLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	   
		
				 VitalSetupHoldCheck (
        Violation      => Tviol_CI_CLK_posedge,
        TimingData     => Tmkr_CI_CLK_posedge,
        TestSignal     => CI_ipd,
        TestSignalName => "CI",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_CI_CLK_posedge_posedge,
        SetupLow       => tsetup_CI_CLK_negedge_posedge,
        HoldLow        => thold_CI_CLK_posedge_posedge,
        HoldHigh       => thold_CI_CLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		
		 VitalSetupHoldCheck (
        Violation      => Tviol_ACCUMCI_CLK_posedge,
        TimingData     => Tmkr_ACCUMCI_CLK_posedge,
        TestSignal     => ACCUMCI_ipd,
        TestSignalName => "ACCUMCI",
        TestDelay      => 0 ns,
        RefSignal      => CLK_ipd,
        RefSignalName  => "CLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_ACCUMCI_CLK_posedge_posedge,
        SetupLow       => tsetup_ACCUMCI_CLK_negedge_posedge,
        HoldLow        => thold_ACCUMCI_CLK_posedge_posedge,
        HoldHigh       => thold_ACCUMCI_CLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
		
		
		 VitalPeriodPulseCheck (
        Violation      => Pviol_CLK,
        PeriodData     => PInfo_CLK,
        TestSignal     => CLK_ipd,
        TestSignalName => "CLK",
        TestDelay      => 0 ns,
        Period         => tperiod_CLK_posedge,
        PulseWidthHigh => tpw_CLK_posedge,
        PulseWidthLow  => tpw_CLK_negedge,
        CheckEnabled   =>true,
        HeaderMsg      => "/SB_MAC16",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
		
		
		VitalRecoveryRemovalCheck (
       Violation               => Tviol_IRSTTOP_CLK_posedge,
       TimingData              => Tmkr_IRSTTOP_CLK_posedge,
       TestSignal              => IRSTTOP_ipd,
       TestSignalName          => "IRSTTOP",
       TestDelay               => 0 ns,
       RefSignal               => CLK_ipd,
       RefSignalName          => "CLK",
       RefDelay                => 0 ns,
       Recovery                => trecovery_IRSTTOP_CLK_negedge_posedge,
       Removal                 => tremoval_IRSTTOP_CLK_negedge_posedge,
       ActiveLow               => FALSE,
       CheckEnabled            => true,
       RefTransition           => 'R',
       HeaderMsg               => "/SB_RAM4KNR",
       Xon                     => Xon,
       MsgOn                   => MsgOn,
       MsgSeverity             => WARNING);
	   
	   VitalRecoveryRemovalCheck (
       Violation               => Tviol_IRSTTOP_CLK_negedge,
       TimingData              => Tmkr_IRSTTOP_CLK_negedge,
       TestSignal              => IRSTTOP_ipd,
       TestSignalName          => "IRSTTOP",
       TestDelay               => 0 ns,
       RefSignal               => CLK_ipd,
       RefSignalName          => "CLK",
       RefDelay                => 0 ns,
       Recovery                => trecovery_IRSTTOP_CLK_posedge_posedge,
       Removal                 => tremoval_IRSTTOP_CLK_posedge_posedge,
       ActiveLow               => FALSE,
       CheckEnabled            => true,
       RefTransition           => 'R',
       HeaderMsg               => "/SB_RAM4KNR",
       Xon                     => Xon,
       MsgOn                   => MsgOn,
       MsgSeverity             => WARNING);
	   
		VitalRecoveryRemovalCheck (
       Violation               => Tviol_IRSTBOT_CLK_negedge,
       TimingData              => Tmkr_IRSTBOT_CLK_negedge,
       TestSignal              => IRSTBOT_ipd,
       TestSignalName          => "IRSTBOT",
       TestDelay               => 0 ns,
       RefSignal               => CLK_ipd,
       RefSignalName          => "CLK",
       RefDelay                => 0 ns,
       Recovery                => trecovery_IRSTBOT_CLK_negedge_posedge,
       Removal                 => tremoval_IRSTBOT_CLK_negedge_posedge,
       ActiveLow               => FALSE,
       CheckEnabled            => true,
       RefTransition           => 'R',
       HeaderMsg               => "/SB_RAM4KNR",
       Xon                     => Xon,
       MsgOn                   => MsgOn,
       MsgSeverity             => WARNING);  

		VitalRecoveryRemovalCheck (
       Violation               => Tviol_IRSTBOT_CLK_posedge,
       TimingData              => Tmkr_IRSTBOT_CLK_posedge,
       TestSignal              => IRSTBOT_ipd,
       TestSignalName          => "IRSTBOT",
       TestDelay               => 0 ns,
       RefSignal               => CLK_ipd,
       RefSignalName          => "CLK",
       RefDelay                => 0 ns,
       Recovery                => trecovery_IRSTBOT_CLK_posedge_posedge,
       Removal                 => tremoval_IRSTBOT_CLK_posedge_posedge,
       ActiveLow               => FALSE,
       CheckEnabled            => true,
       RefTransition           => 'R',
       HeaderMsg               => "/SB_RAM4KNR",
       Xon                     => Xon,
       MsgOn                   => MsgOn,
       MsgSeverity             => WARNING); 	   
	   
	   	VitalRecoveryRemovalCheck (
       Violation               => Tviol_ORSTTOP_CLK_negedge,
       TimingData              => Tmkr_ORSTTOP_CLK_negedge,
       TestSignal              => ORSTTOP_ipd,
       TestSignalName          => "ORSTTOP",
       TestDelay               => 0 ns,
       RefSignal               => CLK_ipd,
       RefSignalName          => "CLK",
       RefDelay                => 0 ns,
       Recovery                => trecovery_ORSTTOP_CLK_negedge_posedge,
       Removal                 => tremoval_ORSTTOP_CLK_negedge_posedge,
       ActiveLow               => FALSE,
       CheckEnabled            => true,
       RefTransition           => 'R',
       HeaderMsg               => "/SB_RAM4KNR",
       Xon                     => Xon,
       MsgOn                   => MsgOn,
       MsgSeverity             => WARNING);  

 	VitalRecoveryRemovalCheck (
       Violation               => Tviol_ORSTTOP_CLK_posedge,
       TimingData              => Tmkr_ORSTTOP_CLK_posedge,
       TestSignal              => ORSTTOP_ipd,
       TestSignalName          => "ORSTTOP",
       TestDelay               => 0 ns,
       RefSignal               => CLK_ipd,
       RefSignalName          => "CLK",
       RefDelay                => 0 ns,
       Recovery                => trecovery_ORSTTOP_CLK_posedge_posedge,
       Removal                 => tremoval_ORSTTOP_CLK_posedge_posedge,
       ActiveLow               => FALSE,
       CheckEnabled            => true,
       RefTransition           => 'R',
       HeaderMsg               => "/SB_RAM4KNR",
       Xon                     => Xon,
       MsgOn                   => MsgOn,
       MsgSeverity             => WARNING);   	   
	   
	   	VitalRecoveryRemovalCheck (
       Violation               => Tviol_ORSTBOT_CLK_negedge,
       TimingData              => Tmkr_ORSTBOT_CLK_negedge,
       TestSignal              => ORSTBOT_ipd,
       TestSignalName          => "ORSTBOT",
       TestDelay               => 0 ns,
       RefSignal               => CLK_ipd,
       RefSignalName          => "CLK",
       RefDelay                => 0 ns,
       Recovery                => trecovery_ORSTBOT_CLK_negedge_posedge,
       Removal                 => tremoval_ORSTBOT_CLK_negedge_posedge,
       ActiveLow               => FALSE,
       CheckEnabled            => true,
       RefTransition           => 'R',
       HeaderMsg               => "/SB_RAM4KNR",
       Xon                     => Xon,
       MsgOn                   => MsgOn,
       MsgSeverity             => WARNING);  

   	VitalRecoveryRemovalCheck (
       Violation               => Tviol_ORSTBOT_CLK_posedge,
       TimingData              => Tmkr_ORSTBOT_CLK_posedge,
       TestSignal              => ORSTBOT_ipd,
       TestSignalName          => "ORSTBOT",
       TestDelay               => 0 ns,
       RefSignal               => CLK_ipd,
       RefSignalName          => "CLK",
       RefDelay                => 0 ns,
       Recovery                => trecovery_ORSTBOT_CLK_posedge_posedge,
       Removal                 => tremoval_ORSTBOT_CLK_posedge_posedge,
       ActiveLow               => FALSE,
       CheckEnabled            => true,
       RefTransition           => 'R',
       HeaderMsg               => "/SB_RAM4KNR",
       Xon                     => Xon,
       MsgOn                   => MsgOn,
       MsgSeverity             => WARNING); 	   
	end if;	
	end process VITALBehavior;
	
	
	VITALPathDelay          : process (Q_zd,QCO_zd,QACCUMCO_zd)
	variable O_GlitchData  : VitalGlitchDataArrayType (31 downto 0); 
	variable CO_GlitchData: VitalGlitchDataType;  
	variable SIGNEXTOUT_GlitchData: VitalGlitchDataType;
	variable ACCUMCO_GlitchData: VitalGlitchDataType;
  	variable O_zd         : std_logic_vector( 31 downto 0);
	variable CO_zd         : std_logic;
	variable ACCUMCO_zd         : std_logic;
	

begin	
	O_zd:=Q_zd ;
	CO_zd := QCO_zd;
	ACCUMCO_zd := QACCUMCO_zd;
      VitalPathDelay01 (
      OutSignal     => O(0),
      GlitchData    => O_GlitchData(0),
      OutSignalName => "O(0)",
      OutTemp       => O_zd(0),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(0), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(0), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(0), true),
						3 => (A_ipd(0)'last_event, tpd_A_O((511 - 31)- 32*15), true),
						4 => (A_ipd(1)'last_event, tpd_A_O((511 - 31)- 32*14), true),
						5 => (A_ipd(2)'last_event, tpd_A_O((511 - 31)- 32*13), true),
						6 => (A_ipd(3)'last_event, tpd_A_O((511 - 31)- 32*12), true),
						7 => (A_ipd(4)'last_event, tpd_A_O((511 - 31)- 32*11), true), 
						8 => (A_ipd(5)'last_event, tpd_A_O((511 - 31)- 32*10), true),
						9 => (A_ipd(6)'last_event, tpd_A_O((511 - 31)- 32*9), true),
						10 => (A_ipd(7)'last_event, tpd_A_O((511 - 31)- 32*8), true),
						11=> (A_ipd(8)'last_event, tpd_A_O((511 - 31)- 32*7), true),
						12 => (A_ipd(9)'last_event, tpd_A_O((511 - 31)- 32*6), true),
						13 => (A_ipd(10)'last_event, tpd_A_O((511 - 31)- 32*5), true),
						14 => (A_ipd(11)'last_event, tpd_A_O((511 - 31)- 32*4), true),
						15 => (A_ipd(12)'last_event, tpd_A_O((511 - 31)- 32*3), true),
						16=> (A_ipd(13)'last_event, tpd_A_O((511 - 31)- 32*2), true),
						17=> (A_ipd(14)'last_event, tpd_A_O((511 - 31)- 32*1), true), 
						18=> (A_ipd(15)'last_event, tpd_A_O((511 - 31)- 32*0), true), 
						19=> (B_ipd(0)'last_event, tpd_B_O((511 - 31)- 32*15), true),
						20 => (B_ipd(1)'last_event, tpd_B_O((511 - 31)- 32*14), true),
						21 => (B_ipd(2)'last_event, tpd_B_O((511 - 31)- 32*13), true),
						22 => (B_ipd(3)'last_event, tpd_B_O((511 - 31)- 32*12), true),
						23=> (B_ipd(4)'last_event, tpd_B_O((511 - 31)- 32*11), true), 
						24=> (B_ipd(5)'last_event, tpd_B_O((511 - 31)- 32*10), true),
						25 => (B_ipd(6)'last_event, tpd_B_O((511 - 31)- 32*9), true),
						26 => (B_ipd(7)'last_event, tpd_B_O((511 - 31)- 32*8), true),
						27=> (B_ipd(8)'last_event, tpd_B_O((511 - 31)- 32*7), true),
						28 => (B_ipd(9)'last_event, tpd_B_O((511 - 31)- 32*6), true),
						29=> (B_ipd(10)'last_event, tpd_B_O((511 - 31)- 32*5), true),
						30 => (B_ipd(11)'last_event, tpd_B_O((511 - 31)- 32*4), true),
						31 => (B_ipd(12)'last_event, tpd_B_O((511 - 31)- 32*3), true),
						32=> (B_ipd(13)'last_event, tpd_B_O((511 - 31)- 32*2), true),
						33=> (B_ipd(14)'last_event, tpd_B_O((511 - 31)- 32*1), true), 
						34=> (B_ipd(15)'last_event, tpd_B_O((511 - 31)- 32*0), true),
						35=> (C_ipd(0)'last_event, tpd_C_O((511 - 31)- 32*15), true),
						36 => (C_ipd(1)'last_event, tpd_C_O((511 - 31)- 32*14), true),
						37 => (C_ipd(2)'last_event, tpd_C_O((511 - 31)- 32*13), true),
						38 => (C_ipd(3)'last_event, tpd_C_O((511 - 31)- 32*12), true),
						39=> (C_ipd(4)'last_event, tpd_C_O((511 - 31)- 32*11), true), 
						40=> (C_ipd(5)'last_event, tpd_C_O((511 - 31)- 32*10), true),
						41 => (C_ipd(6)'last_event, tpd_C_O((511 - 31)- 32*9), true),
						42 => (C_ipd(7)'last_event, tpd_C_O((511 - 31)- 32*8), true),
						43=> (C_ipd(8)'last_event, tpd_C_O((511 - 31)- 32*7), true),
						44 => (C_ipd(9)'last_event, tpd_C_O((511 - 31)- 32*6), true),
						45=> (C_ipd(10)'last_event, tpd_C_O((511 - 31)- 32*5), true),
						46 => (C_ipd(11)'last_event, tpd_C_O((511 - 31)- 32*4), true),
						47 => (C_ipd(12)'last_event, tpd_C_O((511 - 31)- 32*3), true),
						48=> (C_ipd(13)'last_event, tpd_C_O((511 - 31)- 32*2), true),
						49=> (C_ipd(14)'last_event, tpd_C_O((511 - 31)- 32*1), true), 
						50=> (C_ipd(15)'last_event, tpd_C_O((511 - 31)- 32*0), true),
						51=> (D_ipd(0)'last_event, tpd_D_O((511 - 31)- 32*15), true),
						52 => (D_ipd(1)'last_event, tpd_D_O((511 - 31)- 32*14), true),
						53 => (D_ipd(2)'last_event, tpd_D_O((511 - 31)- 32*13), true),
						54 => (D_ipd(3)'last_event, tpd_D_O((511 - 31)- 32*12), true),
						55=> (D_ipd(4)'last_event, tpd_D_O((511 - 31)- 32*11), true), 
						56=> (D_ipd(5)'last_event, tpd_D_O((511 - 31)- 32*10), true),
						57 => (D_ipd(6)'last_event, tpd_D_O((511 - 31)- 32*9), true),
						58 => (D_ipd(7)'last_event, tpd_D_O((511 - 31)- 32*8), true),
						59=> (D_ipd(8)'last_event, tpd_D_O((511 - 31)- 32*7), true),
						60 => (D_ipd(9)'last_event, tpd_D_O((511 - 31)- 32*6), true),
						61=> (D_ipd(10)'last_event, tpd_D_O((511 - 31)- 32*5), true),
						62 => (D_ipd(11)'last_event, tpd_D_O((511 - 31)- 32*4), true),
						63 => (D_ipd(12)'last_event, tpd_D_O((511 - 31)- 32*3), true),
						64=> (D_ipd(13)'last_event, tpd_D_O((511 - 31)- 32*2), true),
						65=> (D_ipd(14)'last_event, tpd_D_O((511 - 31)- 32*1), true), 
						66=> (D_ipd(15)'last_event, tpd_D_O((511 - 31)- 32*0), true),
						67=> (CI_ipd'last_event, tpd_CI_O(0), true),  
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(0), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(0),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(0),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(0),true)
						),  
		Mode          => VitalTransport, 
	 	IgnoreDefaultDelay => TRUE, 
		 RejectFastPath=>TRUE,
     	 Xon           => Xon,
     	 MsgOn         => MsgOn,
     	 MsgSeverity   => warning);	
	  
	  
	  VitalPathDelay01 (
      OutSignal     => O(1),
      GlitchData    => O_GlitchData(1),
      OutSignalName => "O(1)",
      OutTemp       => O_zd(1),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(1), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(1), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(1), true),
						3 => (A_ipd(0)'last_event,  tpd_A_O((511 - 30)- 32*15 ), true),
						4 => (A_ipd(1)'last_event,  tpd_A_O((511 - 30)- 32*14 ), true),
						5 => (A_ipd(2)'last_event,  tpd_A_O((511 - 30)- 32*13 ), true),
						6 => (A_ipd(3)'last_event,  tpd_A_O((511 - 30)- 32*12 ), true),
						7 => (A_ipd(4)'last_event,  tpd_A_O((511 - 30)- 32*11 ), true), 
						8 => (A_ipd(5)'last_event,  tpd_A_O((511 - 30)- 32*10 ), true),
						9 => (A_ipd(6)'last_event,  tpd_A_O((511 - 30)- 32*9 ), true),
						10 => (A_ipd(7)'last_event,  tpd_A_O((511 - 30)- 32*8 ), true),
						11=> (A_ipd(8)'last_event,  tpd_A_O((511 - 30)- 32*7 ), true),
						12 => (A_ipd(9)'last_event,  tpd_A_O((511 - 30)- 32*6 ), true),
						13 => (A_ipd(10)'last_event,  tpd_A_O((511 - 30)- 32*5 ), true),
						14 => (A_ipd(11)'last_event,  tpd_A_O((511 - 30)- 32*4 ), true),
						15 => (A_ipd(12)'last_event,  tpd_A_O((511 - 30)- 32*3 ), true),
						16=> (A_ipd(13)'last_event,  tpd_A_O((511 - 30)- 32*2), true),
						17=> (A_ipd(14)'last_event,  tpd_A_O((511 - 30)- 32*1 ), true), 
						18=> (A_ipd(15)'last_event,  tpd_A_O((511 - 30)- 32*0 ), true), 
						19=> (B_ipd(0)'last_event,  tpd_B_O((511 - 30)- 32*15 ), true),
						20 => (B_ipd(1)'last_event,  tpd_B_O((511 - 30)- 32*14 ), true),
						21 => (B_ipd(2)'last_event,  tpd_B_O((511 - 30)- 32*13 ), true),
						22 => (B_ipd(3)'last_event,  tpd_B_O((511 - 30)- 32*12 ), true),
						23=> (B_ipd(4)'last_event,  tpd_B_O((511 - 30)- 32*11 ), true), 
						24=> (B_ipd(5)'last_event,  tpd_B_O((511 - 30)- 32*10 ), true),
						25 => (B_ipd(6)'last_event,  tpd_B_O((511 - 30)- 32*9 ), true),
						26 => (B_ipd(7)'last_event,  tpd_B_O((511 - 30)- 32*8 ), true),
						27=> (B_ipd(8)'last_event,  tpd_B_O((511 - 30)- 32*7), true),
						28 => (B_ipd(9)'last_event,  tpd_B_O((511 - 30)- 32*6 ), true),
						29=> (B_ipd(10)'last_event,  tpd_B_O((511 - 30)- 32*5 ), true),
						30 => (B_ipd(11)'last_event,  tpd_B_O((511 - 30)- 32*4 ), true),
						31 => (B_ipd(12)'last_event,  tpd_B_O((511 - 30)- 32*3 ), true),
						32=> (B_ipd(13)'last_event,  tpd_B_O((511 - 30)- 32*2 ), true),
						33=> (B_ipd(14)'last_event,  tpd_B_O((511 - 30)- 32*1 ), true), 
						34=> (B_ipd(15)'last_event,  tpd_B_O((511 - 30)- 32*0 ), true),
						35=> (C_ipd(0)'last_event,  tpd_C_O((511 - 30)- 32*15 ), true),
						36 => (C_ipd(1)'last_event,  tpd_C_O((511 - 30)- 32*14 ), true),
						37 => (C_ipd(2)'last_event,  tpd_C_O((511 - 30)- 32*13 ), true),
						38 => (C_ipd(3)'last_event,  tpd_C_O((511 - 30)- 32*12 ), true),
						39=> (C_ipd(4)'last_event,  tpd_C_O((511 - 30)- 32*11 ), true), 
						40=> (C_ipd(5)'last_event,  tpd_C_O((511 - 30)- 32*10 ), true),
						41 => (C_ipd(6)'last_event,  tpd_C_O((511 - 30)- 32*9 ), true),
						42 => (C_ipd(7)'last_event,  tpd_C_O((511 - 30)- 32*8 ), true),
						43=> (C_ipd(8)'last_event,  tpd_C_O((511 - 30)- 32*7), true),
						44 => (C_ipd(9)'last_event,  tpd_C_O((511 - 30)- 32*6 ), true),
						45=> (C_ipd(10)'last_event,  tpd_C_O((511 - 30)- 32*5 ), true),
						46 => (C_ipd(11)'last_event,  tpd_C_O((511 - 30)- 32*4 ), true),
						47 => (C_ipd(12)'last_event,  tpd_C_O((511 - 30)- 32*3 ), true),
						48=> (C_ipd(13)'last_event,  tpd_C_O((511 - 30)- 32*2 ), true),
						49=> (C_ipd(14)'last_event,  tpd_C_O((511 - 30)- 32*1 ), true), 
						50=> (C_ipd(15)'last_event,  tpd_C_O((511 - 30)- 32*0 ), true),
						51=> (D_ipd(0)'last_event,  tpd_D_O((511 - 30)- 32*15 ), true),
						52 => (D_ipd(1)'last_event,  tpd_D_O((511 - 30)- 32*14 ), true),
						53 => (D_ipd(2)'last_event,  tpd_D_O((511 - 30)- 32*13 ), true),
						54 => (D_ipd(3)'last_event,  tpd_D_O((511 - 30)- 32*12 ), true),
						55=> (D_ipd(4)'last_event,  tpd_D_O((511 - 30)- 32*11 ), true), 
						56=> (D_ipd(5)'last_event,  tpd_D_O((511 - 30)- 32*10 ), true),
						57 => (D_ipd(6)'last_event,  tpd_D_O((511 - 30)- 32*9 ), true),
						58 => (D_ipd(7)'last_event,  tpd_D_O((511 - 30)- 32*8 ), true),
						59=> (D_ipd(8)'last_event,  tpd_D_O((511 - 30)- 32*7 ), true),
						60 => (D_ipd(9)'last_event,  tpd_D_O((511 - 30)- 32*6 ), true),
						61=> (D_ipd(10)'last_event,  tpd_D_O((511 - 30)- 32*5 ), true),
						62 => (D_ipd(11)'last_event,  tpd_D_O((511 - 30)- 32*4 ), true),
						63 => (D_ipd(12)'last_event,  tpd_D_O((511 - 30)- 32*3 ), true),
						64=> (D_ipd(13)'last_event,  tpd_D_O((511 - 30)- 32*2 ), true),
						65=> (D_ipd(14)'last_event,  tpd_D_O((511 - 30)- 32*1 ), true), 
						66=> (D_ipd(15)'last_event,  tpd_D_O((511 - 30)- 32*0 ), true),
						67=> (CI_ipd'last_event, tpd_CI_O(1), true),
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(1), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(1),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(1),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(1),true)),
      Mode          => VitalTransport, 
	  IgnoreDefaultDelay => TRUE,
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);	
	  
	  
	    
	  VitalPathDelay01 (
      OutSignal     => O(2),
      GlitchData    => O_GlitchData(2),
      OutSignalName => "O(2)",
      OutTemp       => O_zd(2),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(2), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(2), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(2), true),
						3 => (A_ipd(0)'last_event,  tpd_A_O((511 - 29)- 32*15 ), true),
						4 => (A_ipd(1)'last_event,  tpd_A_O((511 - 29)- 32*14 ), true),
						5 => (A_ipd(2)'last_event,  tpd_A_O((511 - 29)- 32*13 ), true),
						6 => (A_ipd(3)'last_event,  tpd_A_O((511 - 29)- 32*12 ), true),
						7 => (A_ipd(4)'last_event,  tpd_A_O((511 - 29)- 32*11 ), true), 
						8 => (A_ipd(5)'last_event,  tpd_A_O((511 - 29)- 32*10 ), true),
						9 => (A_ipd(6)'last_event,  tpd_A_O((511 - 29)- 32*9 ), true),
						10 => (A_ipd(7)'last_event,  tpd_A_O((511 - 29)- 32*8 ), true),
						11=> (A_ipd(8)'last_event,  tpd_A_O((511 - 29)- 32*7 ), true),
						12 => (A_ipd(9)'last_event,  tpd_A_O((511 - 29)- 32*6 ), true),
						13 => (A_ipd(10)'last_event,  tpd_A_O((511 - 29)- 32*5 ), true),
						14 => (A_ipd(11)'last_event,  tpd_A_O((511 - 29)- 32*4 ), true),
						15 => (A_ipd(12)'last_event,  tpd_A_O((511 - 29)- 32*3 ), true),
						16=> (A_ipd(13)'last_event,  tpd_A_O((511 - 29)- 32*2), true),
						17=> (A_ipd(14)'last_event,  tpd_A_O((511 - 29)- 32*1 ), true), 
						18=> (A_ipd(15)'last_event,  tpd_A_O((511 - 29)- 32*0 ), true), 
						19=> (B_ipd(0)'last_event,  tpd_B_O((511 - 29)- 32*15 ), true),
						20 => (B_ipd(1)'last_event,  tpd_B_O((511 - 29)- 32*14 ), true),
						21 => (B_ipd(2)'last_event,  tpd_B_O((511 - 29)- 32*13 ), true),
						22 => (B_ipd(3)'last_event,  tpd_B_O((511 - 29)- 32*12 ), true),
						23=> (B_ipd(4)'last_event,  tpd_B_O((511 - 29)- 32*11 ), true), 
						24=> (B_ipd(5)'last_event,  tpd_B_O((511 - 29)- 32*10 ), true),
						25 => (B_ipd(6)'last_event,  tpd_B_O((511 - 29)- 32*9 ), true),
						26 => (B_ipd(7)'last_event,  tpd_B_O((511 - 29)- 32*8 ), true),
						27=> (B_ipd(8)'last_event,  tpd_B_O((511 - 29)- 32*7), true),
						28 => (B_ipd(9)'last_event,  tpd_B_O((511 - 29)- 32*6 ), true),
						29=> (B_ipd(10)'last_event,  tpd_B_O((511 - 29)- 32*5 ), true),
						30 => (B_ipd(11)'last_event,  tpd_B_O((511 - 29)- 32*4 ), true),
						31 => (B_ipd(12)'last_event,  tpd_B_O((511 - 29)- 32*3 ), true),
						32=> (B_ipd(13)'last_event,  tpd_B_O((511 - 29)- 32*2 ), true),
						33=> (B_ipd(14)'last_event,  tpd_B_O((511 - 29)- 32*1 ), true), 
						34=> (B_ipd(15)'last_event,  tpd_B_O((511 - 29)- 32*0 ), true),
						35=> (C_ipd(0)'last_event,  tpd_C_O((511 - 29)- 32*15 ), true),
						36 => (C_ipd(1)'last_event,  tpd_C_O((511 - 29)- 32*14 ), true),
						37 => (C_ipd(2)'last_event,  tpd_C_O((511 - 29)- 32*13 ), true),
						38 => (C_ipd(3)'last_event,  tpd_C_O((511 - 29)- 32*12 ), true),
						39=> (C_ipd(4)'last_event,  tpd_C_O((511 - 29)- 32*11 ), true), 
						40=> (C_ipd(5)'last_event,  tpd_C_O((511 - 29)- 32*10 ), true),
						41 => (C_ipd(6)'last_event,  tpd_C_O((511 - 29)- 32*9 ), true),
						42 => (C_ipd(7)'last_event,  tpd_C_O((511 - 29)- 32*8 ), true),
						43=> (C_ipd(8)'last_event,  tpd_C_O((511 - 29)- 32*7), true),
						44 => (C_ipd(9)'last_event,  tpd_C_O((511 - 29)- 32*6 ), true),
						45=> (C_ipd(10)'last_event,  tpd_C_O((511 - 29)- 32*5 ), true),
						46 => (C_ipd(11)'last_event,  tpd_C_O((511 - 29)- 32*4 ), true),
						47 => (C_ipd(12)'last_event,  tpd_C_O((511 - 29)- 32*3 ), true),
						48=> (C_ipd(13)'last_event,  tpd_C_O((511 - 29)- 32*2 ), true),
						49=> (C_ipd(14)'last_event,  tpd_C_O((511 - 29)- 32*1 ), true), 
						50=> (C_ipd(15)'last_event,  tpd_C_O((511 - 29)- 32*0 ), true),
						51=> (D_ipd(0)'last_event,  tpd_D_O((511 - 29)- 32*15 ), true),
						52 => (D_ipd(1)'last_event,  tpd_D_O((511 - 29)- 32*14 ), true),
						53 => (D_ipd(2)'last_event,  tpd_D_O((511 - 29)- 32*13 ), true),
						54 => (D_ipd(3)'last_event,  tpd_D_O((511 - 29)- 32*12 ), true),
						55=> (D_ipd(4)'last_event,  tpd_D_O((511 - 29)- 32*11 ), true), 
						56=> (D_ipd(5)'last_event,  tpd_D_O((511 - 29)- 32*10 ), true),
						57 => (D_ipd(6)'last_event,  tpd_D_O((511 - 29)- 32*9 ), true),
						58 => (D_ipd(7)'last_event,  tpd_D_O((511 - 29)- 32*8 ), true),
						59=> (D_ipd(8)'last_event,  tpd_D_O((511 - 29)- 32*7 ), true),
						60 => (D_ipd(9)'last_event,  tpd_D_O((511 - 29)- 32*6 ), true),
						61=> (D_ipd(10)'last_event,  tpd_D_O((511 - 29)- 32*5 ), true),
						62 => (D_ipd(11)'last_event,  tpd_D_O((511 - 29)- 32*4 ), true),
						63 => (D_ipd(12)'last_event,  tpd_D_O((511 - 29)- 32*3 ), true),
						64=> (D_ipd(13)'last_event,  tpd_D_O((511 - 29)- 32*2 ), true),
						65=> (D_ipd(14)'last_event,  tpd_D_O((511 - 29)- 32*1 ), true), 
						66=> (D_ipd(15)'last_event,  tpd_D_O((511 - 29)- 32*0 ), true),
						67=> (CI_ipd'last_event, tpd_CI_O(2), true)  ,  
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(2), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(2),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(2),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(2),true)),
      Mode          => VitalTransport,
	  IgnoreDefaultDelay => TRUE,
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);			 
	  
	  	  VitalPathDelay01 (
      OutSignal     => O(3),
      GlitchData    => O_GlitchData(3),
      OutSignalName => "O(3)",
      OutTemp       => O_zd(3),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(3), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(3), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(3), true),
						3 => (A_ipd(0)'last_event,  tpd_A_O((511 - 28)- 32*15 ), true),
						4 => (A_ipd(1)'last_event,  tpd_A_O((511 - 28)- 32*14 ), true),
						5 => (A_ipd(2)'last_event,  tpd_A_O((511 - 28)- 32*13 ), true),
						6 => (A_ipd(3)'last_event,  tpd_A_O((511 - 28)- 32*12 ), true),
						7 => (A_ipd(4)'last_event,  tpd_A_O((511 - 28)- 32*11 ), true), 
						8 => (A_ipd(5)'last_event,  tpd_A_O((511 - 28)- 32*10 ), true),
						9 => (A_ipd(6)'last_event,  tpd_A_O((511 - 28)- 32*9 ), true),
						10 => (A_ipd(7)'last_event,  tpd_A_O((511 - 28)- 32*8 ), true),
						11=> (A_ipd(8)'last_event,  tpd_A_O((511 - 28)- 32*7 ), true),
						12 => (A_ipd(9)'last_event,  tpd_A_O((511 - 28)- 32*6 ), true),
						13 => (A_ipd(10)'last_event,  tpd_A_O((511 - 28)- 32*5 ), true),
						14 => (A_ipd(11)'last_event,  tpd_A_O((511 - 28)- 32*4 ), true),
						15 => (A_ipd(12)'last_event,  tpd_A_O((511 - 28)- 32*3 ), true),
						16=> (A_ipd(13)'last_event,  tpd_A_O((511 - 28)- 32*2), true),
						17=> (A_ipd(14)'last_event,  tpd_A_O((511 - 28)- 32*1 ), true), 
						18=> (A_ipd(15)'last_event,  tpd_A_O((511 - 28)- 32*0 ), true), 
						19=> (B_ipd(0)'last_event,  tpd_B_O((511 - 28)- 32*15 ), true),
						20 => (B_ipd(1)'last_event,  tpd_B_O((511 - 28)- 32*14 ), true),
						21 => (B_ipd(2)'last_event,  tpd_B_O((511 - 28)- 32*13 ), true),
						22 => (B_ipd(3)'last_event,  tpd_B_O((511 - 28)- 32*12 ), true),
						23=> (B_ipd(4)'last_event,  tpd_B_O((511 - 28)- 32*11 ), true), 
						24=> (B_ipd(5)'last_event,  tpd_B_O((511 - 28)- 32*10 ), true),
						25 => (B_ipd(6)'last_event,  tpd_B_O((511 - 28)- 32*9 ), true),
						26 => (B_ipd(7)'last_event,  tpd_B_O((511 - 28)- 32*8 ), true),
						27=> (B_ipd(8)'last_event,  tpd_B_O((511 - 28)- 32*7), true),
						28 => (B_ipd(9)'last_event,  tpd_B_O((511 - 28)- 32*6 ), true),
						29=> (B_ipd(10)'last_event,  tpd_B_O((511 - 28)- 32*5 ), true),
						30 => (B_ipd(11)'last_event,  tpd_B_O((511 - 28)- 32*4 ), true),
						31 => (B_ipd(12)'last_event,  tpd_B_O((511 - 28)- 32*3 ), true),
						32=> (B_ipd(13)'last_event,  tpd_B_O((511 - 28)- 32*2 ), true),
						33=> (B_ipd(14)'last_event,  tpd_B_O((511 - 28)- 32*1 ), true), 
						34=> (B_ipd(15)'last_event,  tpd_B_O((511 - 28)- 32*0 ), true),
						35=> (C_ipd(0)'last_event,  tpd_C_O((511 - 28)- 32*15 ), true),
						36 => (C_ipd(1)'last_event,  tpd_C_O((511 - 28)- 32*14 ), true),
						37 => (C_ipd(2)'last_event,  tpd_C_O((511 - 28)- 32*13 ), true),
						38 => (C_ipd(3)'last_event,  tpd_C_O((511 - 28)- 32*12 ), true),
						39=> (C_ipd(4)'last_event,  tpd_C_O((511 - 28)- 32*11 ), true), 
						40=> (C_ipd(5)'last_event,  tpd_C_O((511 - 28)- 32*10 ), true),
						41 => (C_ipd(6)'last_event,  tpd_C_O((511 - 28)- 32*9 ), true),
						42 => (C_ipd(7)'last_event,  tpd_C_O((511 - 28)- 32*8 ), true),
						43=> (C_ipd(8)'last_event,  tpd_C_O((511 - 28)- 32*7), true),
						44 => (C_ipd(9)'last_event,  tpd_C_O((511 - 28)- 32*6 ), true),
						45=> (C_ipd(10)'last_event,  tpd_C_O((511 - 28)- 32*5 ), true),
						46 => (C_ipd(11)'last_event,  tpd_C_O((511 - 28)- 32*4 ), true),
						47 => (C_ipd(12)'last_event,  tpd_C_O((511 - 28)- 32*3 ), true),
						48=> (C_ipd(13)'last_event,  tpd_C_O((511 - 28)- 32*2 ), true),
						49=> (C_ipd(14)'last_event,  tpd_C_O((511 - 28)- 32*1 ), true), 
						50=> (C_ipd(15)'last_event,  tpd_C_O((511 - 28)- 32*0 ), true),
						51=> (D_ipd(0)'last_event,  tpd_D_O((511 - 28)- 32*15 ), true),
						52 => (D_ipd(1)'last_event,  tpd_D_O((511 - 28)- 32*14 ), true),
						53 => (D_ipd(2)'last_event,  tpd_D_O((511 - 28)- 32*13 ), true),
						54 => (D_ipd(3)'last_event,  tpd_D_O((511 - 28)- 32*12 ), true),
						55=> (D_ipd(4)'last_event,  tpd_D_O((511 - 28)- 32*11 ), true), 
						56=> (D_ipd(5)'last_event,  tpd_D_O((511 - 28)- 32*10 ), true),
						57 => (D_ipd(6)'last_event,  tpd_D_O((511 - 28)- 32*9 ), true),
						58 => (D_ipd(7)'last_event,  tpd_D_O((511 - 28)- 32*8 ), true),
						59=> (D_ipd(8)'last_event,  tpd_D_O((511 - 28)- 32*7 ), true),
						60 => (D_ipd(9)'last_event,  tpd_D_O((511 - 28)- 32*6 ), true),
						61=> (D_ipd(10)'last_event,  tpd_D_O((511 - 28)- 32*5 ), true),
						62 => (D_ipd(11)'last_event,  tpd_D_O((511 - 28)- 32*4 ), true),
						63 => (D_ipd(12)'last_event,  tpd_D_O((511 - 28)- 32*3 ), true),
						64=> (D_ipd(13)'last_event,  tpd_D_O((511 - 28)- 32*2 ), true),
						65=> (D_ipd(14)'last_event,  tpd_D_O((511 - 28)- 32*1 ), true), 
						66=> (D_ipd(15)'last_event,  tpd_D_O((511 - 28)- 32*0 ), true),
						67=> (CI_ipd'last_event, tpd_CI_O(3), true)  ,  
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(3), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(3),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(3),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(3),true)),
      Mode          => VitalTransport,
	  IgnoreDefaultDelay => TRUE,
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);	
	      
	  VitalPathDelay01 (
      OutSignal     => O(4),
      GlitchData    => O_GlitchData(4),
      OutSignalName => "O(4)",
      OutTemp       => O_zd(4),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(4), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(4), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(4), true),
						3 => (A_ipd(0)'last_event,  tpd_A_O((511 - 27)- 32*15 ), true),
						4 => (A_ipd(1)'last_event,  tpd_A_O((511 - 27)- 32*14 ), true),
						5 => (A_ipd(2)'last_event,  tpd_A_O((511 - 27)- 32*13 ), true),
						6 => (A_ipd(3)'last_event,  tpd_A_O((511 - 27)- 32*12 ), true),
						7 => (A_ipd(4)'last_event,  tpd_A_O((511 - 27)- 32*11 ), true), 
						8 => (A_ipd(5)'last_event,  tpd_A_O((511 - 27)- 32*10 ), true),
						9 => (A_ipd(6)'last_event,  tpd_A_O((511 - 27)- 32*9 ), true),
						10 => (A_ipd(7)'last_event,  tpd_A_O((511 - 27)- 32*8 ), true),
						11=> (A_ipd(8)'last_event,  tpd_A_O((511 - 27)- 32*7 ), true),
						12 => (A_ipd(9)'last_event,  tpd_A_O((511 - 27)- 32*6 ), true),
						13 => (A_ipd(10)'last_event,  tpd_A_O((511 - 27)- 32*5 ), true),
						14 => (A_ipd(11)'last_event,  tpd_A_O((511 - 27)- 32*4 ), true),
						15 => (A_ipd(12)'last_event,  tpd_A_O((511 - 27)- 32*3 ), true),
						16=> (A_ipd(13)'last_event,  tpd_A_O((511 - 27)- 32*2), true),
						17=> (A_ipd(14)'last_event,  tpd_A_O((511 - 27)- 32*1 ), true), 
						18=> (A_ipd(15)'last_event,  tpd_A_O((511 - 27)- 32*0 ), true), 
						19=> (B_ipd(0)'last_event,  tpd_B_O((511 - 27)- 32*15 ), true),
						20 => (B_ipd(1)'last_event,  tpd_B_O((511 - 27)- 32*14 ), true),
						21 => (B_ipd(2)'last_event,  tpd_B_O((511 - 27)- 32*13 ), true),
						22 => (B_ipd(3)'last_event,  tpd_B_O((511 - 27)- 32*12 ), true),
						23=> (B_ipd(4)'last_event,  tpd_B_O((511 - 27)- 32*11 ), true), 
						24=> (B_ipd(5)'last_event,  tpd_B_O((511 - 27)- 32*10 ), true),
						25 => (B_ipd(6)'last_event,  tpd_B_O((511 - 27)- 32*9 ), true),
						26 => (B_ipd(7)'last_event,  tpd_B_O((511 - 27)- 32*8 ), true),
						27=> (B_ipd(8)'last_event,  tpd_B_O((511 - 27)- 32*7), true),
						28 => (B_ipd(9)'last_event,  tpd_B_O((511 - 27)- 32*6 ), true),
						29=> (B_ipd(10)'last_event,  tpd_B_O((511 - 27)- 32*5 ), true),
						30 => (B_ipd(11)'last_event,  tpd_B_O((511 - 27)- 32*4 ), true),
						31 => (B_ipd(12)'last_event,  tpd_B_O((511 - 27)- 32*3 ), true),
						32=> (B_ipd(13)'last_event,  tpd_B_O((511 - 27)- 32*2 ), true),
						33=> (B_ipd(14)'last_event,  tpd_B_O((511 - 27)- 32*1 ), true), 
						34=> (B_ipd(15)'last_event,  tpd_B_O((511 - 27)- 32*0 ), true),
						35=> (C_ipd(0)'last_event,  tpd_C_O((511 - 27)- 32*15 ), true),
						36 => (C_ipd(1)'last_event,  tpd_C_O((511 - 27)- 32*14 ), true),
						37 => (C_ipd(2)'last_event,  tpd_C_O((511 - 27)- 32*13 ), true),
						38 => (C_ipd(3)'last_event,  tpd_C_O((511 - 27)- 32*12 ), true),
						39=> (C_ipd(4)'last_event,  tpd_C_O((511 - 27)- 32*11 ), true), 
						40=> (C_ipd(5)'last_event,  tpd_C_O((511 - 27)- 32*10 ), true),
						41 => (C_ipd(6)'last_event,  tpd_C_O((511 - 27)- 32*9 ), true),
						42 => (C_ipd(7)'last_event,  tpd_C_O((511 - 27)- 32*8 ), true),
						43=> (C_ipd(8)'last_event,  tpd_C_O((511 - 27)- 32*7), true),
						44 => (C_ipd(9)'last_event,  tpd_C_O((511 - 27)- 32*6 ), true),
						45=> (C_ipd(10)'last_event,  tpd_C_O((511 - 27)- 32*5 ), true),
						46 => (C_ipd(11)'last_event,  tpd_C_O((511 - 27)- 32*4 ), true),
						47 => (C_ipd(12)'last_event,  tpd_C_O((511 - 27)- 32*3 ), true),
						48=> (C_ipd(13)'last_event,  tpd_C_O((511 - 27)- 32*2 ), true),
						49=> (C_ipd(14)'last_event,  tpd_C_O((511 - 27)- 32*1 ), true), 
						50=> (C_ipd(15)'last_event,  tpd_C_O((511 - 27)- 32*0 ), true),
						51=> (D_ipd(0)'last_event,  tpd_D_O((511 - 27)- 32*15 ), true),
						52 => (D_ipd(1)'last_event,  tpd_D_O((511 - 27)- 32*14 ), true),
						53 => (D_ipd(2)'last_event,  tpd_D_O((511 - 27)- 32*13 ), true),
						54 => (D_ipd(3)'last_event,  tpd_D_O((511 - 27)- 32*12 ), true),
						55=> (D_ipd(4)'last_event,  tpd_D_O((511 - 27)- 32*11 ), true), 
						56=> (D_ipd(5)'last_event,  tpd_D_O((511 - 27)- 32*10 ), true),
						57 => (D_ipd(6)'last_event,  tpd_D_O((511 - 27)- 32*9 ), true),
						58 => (D_ipd(7)'last_event,  tpd_D_O((511 - 27)- 32*8 ), true),
						59=> (D_ipd(8)'last_event,  tpd_D_O((511 - 27)- 32*7 ), true),
						60 => (D_ipd(9)'last_event,  tpd_D_O((511 - 27)- 32*6 ), true),
						61=> (D_ipd(10)'last_event,  tpd_D_O((511 - 27)- 32*5 ), true),
						62 => (D_ipd(11)'last_event,  tpd_D_O((511 - 27)- 32*4 ), true),
						63 => (D_ipd(12)'last_event,  tpd_D_O((511 - 27)- 32*3 ), true),
						64=> (D_ipd(13)'last_event,  tpd_D_O((511 - 27)- 32*2 ), true),
						65=> (D_ipd(14)'last_event,  tpd_D_O((511 - 27)- 32*1 ), true), 
						66=> (D_ipd(15)'last_event,  tpd_D_O((511 - 27)- 32*0 ), true),
						67=> (CI_ipd'last_event, tpd_CI_O(4), true)  ,  
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(4), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(4),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(4),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(4),true)),
      Mode          => VitalTransport,	  
	  IgnoreDefaultDelay => TRUE, 
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);
	  
	      

	  
	  
	      
	  VitalPathDelay01 (
      OutSignal     => O(5),
      GlitchData    => O_GlitchData(5),
      OutSignalName => "O(5)",
      OutTemp       => O_zd(5),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(5), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(5), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(5), true),
						3 => (A_ipd(0)'last_event,  tpd_A_O((511 - 26)- 32*15 ), true),
						4 => (A_ipd(1)'last_event,  tpd_A_O((511 - 26)- 32*14 ), true),
						5 => (A_ipd(2)'last_event,  tpd_A_O((511 - 26)- 32*13 ), true),
						6 => (A_ipd(3)'last_event,  tpd_A_O((511 - 26)- 32*12 ), true),
						7 => (A_ipd(4)'last_event,  tpd_A_O((511 - 26)- 32*11 ), true), 
						8 => (A_ipd(5)'last_event,  tpd_A_O((511 - 26)- 32*10 ), true),
						9 => (A_ipd(6)'last_event,  tpd_A_O((511 - 26)- 32*9 ), true),
						10 => (A_ipd(7)'last_event,  tpd_A_O((511 - 26)- 32*8 ), true),
						11=> (A_ipd(8)'last_event,  tpd_A_O((511 - 26)- 32*7 ), true),
						12 => (A_ipd(9)'last_event,  tpd_A_O((511 - 26)- 32*6 ), true),
						13 => (A_ipd(10)'last_event,  tpd_A_O((511 - 26)- 32*5 ), true),
						14 => (A_ipd(11)'last_event,  tpd_A_O((511 - 26)- 32*4 ), true),
						15 => (A_ipd(12)'last_event,  tpd_A_O((511 - 26)- 32*3 ), true),
						16=> (A_ipd(13)'last_event,  tpd_A_O((511 - 26)- 32*2), true),
						17=> (A_ipd(14)'last_event,  tpd_A_O((511 - 26)- 32*1 ), true), 
						18=> (A_ipd(15)'last_event,  tpd_A_O((511 - 26)- 32*0 ), true), 
						19=> (B_ipd(0)'last_event,  tpd_B_O((511 - 26)- 32*15 ), true),
						20 => (B_ipd(1)'last_event,  tpd_B_O((511 - 26)- 32*14 ), true),
						21 => (B_ipd(2)'last_event,  tpd_B_O((511 - 26)- 32*13 ), true),
						22 => (B_ipd(3)'last_event,  tpd_B_O((511 - 26)- 32*12 ), true),
						23=> (B_ipd(4)'last_event,  tpd_B_O((511 - 26)- 32*11 ), true), 
						24=> (B_ipd(5)'last_event,  tpd_B_O((511 - 26)- 32*10 ), true),
						25 => (B_ipd(6)'last_event,  tpd_B_O((511 - 26)- 32*9 ), true),
						26 => (B_ipd(7)'last_event,  tpd_B_O((511 - 26)- 32*8 ), true),
						27=> (B_ipd(8)'last_event,  tpd_B_O((511 - 26)- 32*7), true),
						28 => (B_ipd(9)'last_event,  tpd_B_O((511 - 26)- 32*6 ), true),
						29=> (B_ipd(10)'last_event,  tpd_B_O((511 - 26)- 32*5 ), true),
						30 => (B_ipd(11)'last_event,  tpd_B_O((511 - 26)- 32*4 ), true),
						31 => (B_ipd(12)'last_event,  tpd_B_O((511 - 26)- 32*3 ), true),
						32=> (B_ipd(13)'last_event,  tpd_B_O((511 - 26)- 32*2 ), true),
						33=> (B_ipd(14)'last_event,  tpd_B_O((511 - 26)- 32*1 ), true), 
						34=> (B_ipd(15)'last_event,  tpd_B_O((511 - 26)- 32*0 ), true),
						35=> (C_ipd(0)'last_event,  tpd_C_O((511 - 26)- 32*15 ), true),
						36 => (C_ipd(1)'last_event,  tpd_C_O((511 - 26)- 32*14 ), true),
						37 => (C_ipd(2)'last_event,  tpd_C_O((511 - 26)- 32*13 ), true),
						38 => (C_ipd(3)'last_event,  tpd_C_O((511 - 26)- 32*12 ), true),
						39=> (C_ipd(4)'last_event,  tpd_C_O((511 - 26)- 32*11 ), true), 
						40=> (C_ipd(5)'last_event,  tpd_C_O((511 - 26)- 32*10 ), true),
						41 => (C_ipd(6)'last_event,  tpd_C_O((511 - 26)- 32*9 ), true),
						42 => (C_ipd(7)'last_event,  tpd_C_O((511 - 26)- 32*8 ), true),
						43=> (C_ipd(8)'last_event,  tpd_C_O((511 - 26)- 32*7), true),
						44 => (C_ipd(9)'last_event,  tpd_C_O((511 - 26)- 32*6 ), true),
						45=> (C_ipd(10)'last_event,  tpd_C_O((511 - 26)- 32*5 ), true),
						46 => (C_ipd(11)'last_event,  tpd_C_O((511 - 26)- 32*4 ), true),
						47 => (C_ipd(12)'last_event,  tpd_C_O((511 - 26)- 32*3 ), true),
						48=> (C_ipd(13)'last_event,  tpd_C_O((511 - 26)- 32*2 ), true),
						49=> (C_ipd(14)'last_event,  tpd_C_O((511 - 26)- 32*1 ), true), 
						50=> (C_ipd(15)'last_event,  tpd_C_O((511 - 26)- 32*0 ), true),
						51=> (D_ipd(0)'last_event,  tpd_D_O((511 - 26)- 32*15 ), true),
						52 => (D_ipd(1)'last_event,  tpd_D_O((511 - 26)- 32*14 ), true),
						53 => (D_ipd(2)'last_event,  tpd_D_O((511 - 26)- 32*13 ), true),
						54 => (D_ipd(3)'last_event,  tpd_D_O((511 - 26)- 32*12 ), true),
						55=> (D_ipd(4)'last_event,  tpd_D_O((511 - 26)- 32*11 ), true), 
						56=> (D_ipd(5)'last_event,  tpd_D_O((511 - 26)- 32*10 ), true),
						57 => (D_ipd(6)'last_event,  tpd_D_O((511 - 26)- 32*9 ), true),
						58 => (D_ipd(7)'last_event,  tpd_D_O((511 - 26)- 32*8 ), true),
						59=> (D_ipd(8)'last_event,  tpd_D_O((511 - 26)- 32*7 ), true),
						60 => (D_ipd(9)'last_event,  tpd_D_O((511 - 26)- 32*6 ), true),
						61=> (D_ipd(10)'last_event,  tpd_D_O((511 - 26)- 32*5 ), true),
						62 => (D_ipd(11)'last_event,  tpd_D_O((511 - 26)- 32*4 ), true),
						63 => (D_ipd(12)'last_event,  tpd_D_O((511 - 26)- 32*3 ), true),
						64=> (D_ipd(13)'last_event,  tpd_D_O((511 - 26)- 32*2 ), true),
						65=> (D_ipd(14)'last_event,  tpd_D_O((511 - 26)- 32*1 ), true), 
						66=> (D_ipd(15)'last_event,  tpd_D_O((511 - 26)- 32*0 ), true),
						67=> (CI_ipd'last_event, tpd_CI_O(5), true)  ,  
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(5), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(5),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(5),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(5),true)),
      Mode          => VitalTransport, 
	  IgnoreDefaultDelay => TRUE,
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);
	  
	   VitalPathDelay01 (
      OutSignal     => O(6),
      GlitchData    => O_GlitchData(6),
      OutSignalName => "O(6)",
      OutTemp       => O_zd(6),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(6), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(6), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(6), true),
							3 => (A_ipd(0)'last_event,  tpd_A_O((511 - 25)- 32*15 ), true),
						4 => (A_ipd(1)'last_event,  tpd_A_O((511 - 25)- 32*14 ), true),
						5 => (A_ipd(2)'last_event,  tpd_A_O((511 - 25)- 32*13 ), true),
						6 => (A_ipd(3)'last_event,  tpd_A_O((511 - 25)- 32*12 ), true),
						7 => (A_ipd(4)'last_event,  tpd_A_O((511 - 25)- 32*11 ), true), 
						8 => (A_ipd(5)'last_event,  tpd_A_O((511 - 25)- 32*10 ), true),
						9 => (A_ipd(6)'last_event,  tpd_A_O((511 - 25)- 32*9 ), true),
						10 => (A_ipd(7)'last_event,  tpd_A_O((511 - 25)- 32*8 ), true),
						11=> (A_ipd(8)'last_event,  tpd_A_O((511 - 25)- 32*7 ), true),
						12 => (A_ipd(9)'last_event,  tpd_A_O((511 - 25)- 32*6 ), true),
						13 => (A_ipd(10)'last_event,  tpd_A_O((511 - 25)- 32*5 ), true),
						14 => (A_ipd(11)'last_event,  tpd_A_O((511 - 25)- 32*4 ), true),
						15 => (A_ipd(12)'last_event,  tpd_A_O((511 - 25)- 32*3 ), true),
						16=> (A_ipd(13)'last_event,  tpd_A_O((511 - 25)- 32*2), true),
						17=> (A_ipd(14)'last_event,  tpd_A_O((511 - 25)- 32*1 ), true), 
						18=> (A_ipd(15)'last_event,  tpd_A_O((511 - 25)- 32*0 ), true), 
						19=> (B_ipd(0)'last_event,  tpd_B_O((511 - 25)- 32*15 ), true),
						20 => (B_ipd(1)'last_event,  tpd_B_O((511 - 25)- 32*14 ), true),
						21 => (B_ipd(2)'last_event,  tpd_B_O((511 - 25)- 32*13 ), true),
						22 => (B_ipd(3)'last_event,  tpd_B_O((511 - 25)- 32*12 ), true),
						23=> (B_ipd(4)'last_event,  tpd_B_O((511 - 25)- 32*11 ), true), 
						24=> (B_ipd(5)'last_event,  tpd_B_O((511 - 25)- 32*10 ), true),
						25 => (B_ipd(6)'last_event,  tpd_B_O((511 - 25)- 32*9 ), true),
						26 => (B_ipd(7)'last_event,  tpd_B_O((511 - 25)- 32*8 ), true),
						27=> (B_ipd(8)'last_event,  tpd_B_O((511 - 25)- 32*7), true),
						28 => (B_ipd(9)'last_event,  tpd_B_O((511 - 25)- 32*6 ), true),
						29=> (B_ipd(10)'last_event,  tpd_B_O((511 - 25)- 32*5 ), true),
						30 => (B_ipd(11)'last_event,  tpd_B_O((511 - 25)- 32*4 ), true),
						31 => (B_ipd(12)'last_event,  tpd_B_O((511 - 25)- 32*3 ), true),
						32=> (B_ipd(13)'last_event,  tpd_B_O((511 - 25)- 32*2 ), true),
						33=> (B_ipd(14)'last_event,  tpd_B_O((511 - 25)- 32*1 ), true), 
						34=> (B_ipd(15)'last_event,  tpd_B_O((511 - 25)- 32*0 ), true),
						35=> (C_ipd(0)'last_event,  tpd_C_O((511 - 25)- 32*15 ), true),
						36 => (C_ipd(1)'last_event,  tpd_C_O((511 - 25)- 32*14 ), true),
						37 => (C_ipd(2)'last_event,  tpd_C_O((511 - 25)- 32*13 ), true),
						38 => (C_ipd(3)'last_event,  tpd_C_O((511 - 25)- 32*12 ), true),
						39=> (C_ipd(4)'last_event,  tpd_C_O((511 - 25)- 32*11 ), true), 
						40=> (C_ipd(5)'last_event,  tpd_C_O((511 - 25)- 32*10 ), true),
						41 => (C_ipd(6)'last_event,  tpd_C_O((511 - 25)- 32*9 ), true),
						42 => (C_ipd(7)'last_event,  tpd_C_O((511 - 25)- 32*8 ), true),
						43=> (C_ipd(8)'last_event,  tpd_C_O((511 - 25)- 32*7), true),
						44 => (C_ipd(9)'last_event,  tpd_C_O((511 - 25)- 32*6 ), true),
						45=> (C_ipd(10)'last_event,  tpd_C_O((511 - 25)- 32*5 ), true),
						46 => (C_ipd(11)'last_event,  tpd_C_O((511 - 25)- 32*4 ), true),
						47 => (C_ipd(12)'last_event,  tpd_C_O((511 - 25)- 32*3 ), true),
						48=> (C_ipd(13)'last_event,  tpd_C_O((511 - 25)- 32*2 ), true),
						49=> (C_ipd(14)'last_event,  tpd_C_O((511 - 25)- 32*1 ), true), 
						50=> (C_ipd(15)'last_event,  tpd_C_O((511 - 25)- 32*0 ), true),
						51=> (D_ipd(0)'last_event,  tpd_D_O((511 - 25)- 32*15 ), true),
						52 => (D_ipd(1)'last_event,  tpd_D_O((511 - 25)- 32*14 ), true),
						53 => (D_ipd(2)'last_event,  tpd_D_O((511 - 25)- 32*13 ), true),
						54 => (D_ipd(3)'last_event,  tpd_D_O((511 - 25)- 32*12 ), true),
						55=> (D_ipd(4)'last_event,  tpd_D_O((511 - 25)- 32*11 ), true), 
						56=> (D_ipd(5)'last_event,  tpd_D_O((511 - 25)- 32*10 ), true),
						57 => (D_ipd(6)'last_event,  tpd_D_O((511 - 25)- 32*9 ), true),
						58 => (D_ipd(7)'last_event,  tpd_D_O((511 - 25)- 32*8 ), true),
						59=> (D_ipd(8)'last_event,  tpd_D_O((511 - 25)- 32*7 ), true),
						60 => (D_ipd(9)'last_event,  tpd_D_O((511 - 25)- 32*6 ), true),
						61=> (D_ipd(10)'last_event,  tpd_D_O((511 - 25)- 32*5 ), true),
						62 => (D_ipd(11)'last_event,  tpd_D_O((511 - 25)- 32*4 ), true),
						63 => (D_ipd(12)'last_event,  tpd_D_O((511 - 25)- 32*3 ), true),
						64=> (D_ipd(13)'last_event,  tpd_D_O((511 - 25)- 32*2 ), true),
						65=> (D_ipd(14)'last_event,  tpd_D_O((511 - 25)- 32*1 ), true), 
						66=> (D_ipd(15)'last_event,  tpd_D_O((511 - 25)- 32*0 ), true),
						67=> (CI_ipd'last_event, tpd_CI_O(6), true)  ,  
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(6), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(6),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(6),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(6),true)),
      Mode          => VitalTransport,	  
	  IgnoreDefaultDelay => TRUE,
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);
	  
	  	   VitalPathDelay01 (
      OutSignal     => O(7),
      GlitchData    => O_GlitchData(7),
      OutSignalName => "O(7)",
      OutTemp       => O_zd(7),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(7), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(7), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(7), true),
							3 => (A_ipd(0)'last_event,  tpd_A_O((511 - 24)- 32*15 ), true),
						4 => (A_ipd(1)'last_event,  tpd_A_O((511 - 24)- 32*14 ), true),
						5 => (A_ipd(2)'last_event,  tpd_A_O((511 - 24)- 32*13 ), true),
						6 => (A_ipd(3)'last_event,  tpd_A_O((511 - 24)- 32*12 ), true),
						7 => (A_ipd(4)'last_event,  tpd_A_O((511 - 24)- 32*11 ), true), 
						8 => (A_ipd(5)'last_event,  tpd_A_O((511 - 24)- 32*10 ), true),
						9 => (A_ipd(6)'last_event,  tpd_A_O((511 - 24)- 32*9 ), true),
						10 => (A_ipd(7)'last_event,  tpd_A_O((511 - 24)- 32*8 ), true),
						11=> (A_ipd(8)'last_event,  tpd_A_O((511 - 24)- 32*7 ), true),
						12 => (A_ipd(9)'last_event,  tpd_A_O((511 - 24)- 32*6 ), true),
						13 => (A_ipd(10)'last_event,  tpd_A_O((511 - 24)- 32*5 ), true),
						14 => (A_ipd(11)'last_event,  tpd_A_O((511 - 24)- 32*4 ), true),
						15 => (A_ipd(12)'last_event,  tpd_A_O((511 - 24)- 32*3 ), true),
						16=> (A_ipd(13)'last_event,  tpd_A_O((511 - 24)- 32*2), true),
						17=> (A_ipd(14)'last_event,  tpd_A_O((511 - 24)- 32*1 ), true), 
						18=> (A_ipd(15)'last_event,  tpd_A_O((511 - 24)- 32*0 ), true), 
						19=> (B_ipd(0)'last_event,  tpd_B_O((511 - 24)- 32*15 ), true),
						20 => (B_ipd(1)'last_event,  tpd_B_O((511 - 24)- 32*14 ), true),
						21 => (B_ipd(2)'last_event,  tpd_B_O((511 - 24)- 32*13 ), true),
						22 => (B_ipd(3)'last_event,  tpd_B_O((511 - 24)- 32*12 ), true),
						23=> (B_ipd(4)'last_event,  tpd_B_O((511 - 24)- 32*11 ), true), 
						24=> (B_ipd(5)'last_event,  tpd_B_O((511 - 24)- 32*10 ), true),
						25 => (B_ipd(6)'last_event,  tpd_B_O((511 - 24)- 32*9 ), true),
						26 => (B_ipd(7)'last_event,  tpd_B_O((511 - 24)- 32*8 ), true),
						27=> (B_ipd(8)'last_event,  tpd_B_O((511 - 24)- 32*7), true),
						28 => (B_ipd(9)'last_event,  tpd_B_O((511 - 24)- 32*6 ), true),
						29=> (B_ipd(10)'last_event,  tpd_B_O((511 - 24)- 32*5 ), true),
						30 => (B_ipd(11)'last_event,  tpd_B_O((511 - 24)- 32*4 ), true),
						31 => (B_ipd(12)'last_event,  tpd_B_O((511 - 24)- 32*3 ), true),
						32=> (B_ipd(13)'last_event,  tpd_B_O((511 - 24)- 32*2 ), true),
						33=> (B_ipd(14)'last_event,  tpd_B_O((511 - 24)- 32*1 ), true), 
						34=> (B_ipd(15)'last_event,  tpd_B_O((511 - 24)- 32*0 ), true),
						35=> (C_ipd(0)'last_event,  tpd_C_O((511 - 24)- 32*15 ), true),
						36 => (C_ipd(1)'last_event,  tpd_C_O((511 - 24)- 32*14 ), true),
						37 => (C_ipd(2)'last_event,  tpd_C_O((511 - 24)- 32*13 ), true),
						38 => (C_ipd(3)'last_event,  tpd_C_O((511 - 24)- 32*12 ), true),
						39=> (C_ipd(4)'last_event,  tpd_C_O((511 - 24)- 32*11 ), true), 
						40=> (C_ipd(5)'last_event,  tpd_C_O((511 - 24)- 32*10 ), true),
						41 => (C_ipd(6)'last_event,  tpd_C_O((511 - 24)- 32*9 ), true),
						42 => (C_ipd(7)'last_event,  tpd_C_O((511 - 24)- 32*8 ), true),
						43=> (C_ipd(8)'last_event,  tpd_C_O((511 - 24)- 32*7), true),
						44 => (C_ipd(9)'last_event,  tpd_C_O((511 - 24)- 32*6 ), true),
						45=> (C_ipd(10)'last_event,  tpd_C_O((511 - 24)- 32*5 ), true),
						46 => (C_ipd(11)'last_event,  tpd_C_O((511 - 24)- 32*4 ), true),
						47 => (C_ipd(12)'last_event,  tpd_C_O((511 - 24)- 32*3 ), true),
						48=> (C_ipd(13)'last_event,  tpd_C_O((511 - 24)- 32*2 ), true),
						49=> (C_ipd(14)'last_event,  tpd_C_O((511 - 24)- 32*1 ), true), 
						50=> (C_ipd(15)'last_event,  tpd_C_O((511 - 24)- 32*0 ), true),
						51=> (D_ipd(0)'last_event,  tpd_D_O((511 - 24)- 32*15 ), true),
						52 => (D_ipd(1)'last_event,  tpd_D_O((511 - 24)- 32*14 ), true),
						53 => (D_ipd(2)'last_event,  tpd_D_O((511 - 24)- 32*13 ), true),
						54 => (D_ipd(3)'last_event,  tpd_D_O((511 - 24)- 32*12 ), true),
						55=> (D_ipd(4)'last_event,  tpd_D_O((511 - 24)- 32*11 ), true), 
						56=> (D_ipd(5)'last_event,  tpd_D_O((511 - 24)- 32*10 ), true),
						57 => (D_ipd(6)'last_event,  tpd_D_O((511 - 24)- 32*9 ), true),
						58 => (D_ipd(7)'last_event,  tpd_D_O((511 - 24)- 32*8 ), true),
						59=> (D_ipd(8)'last_event,  tpd_D_O((511 - 24)- 32*7 ), true),
						60 => (D_ipd(9)'last_event,  tpd_D_O((511 - 24)- 32*6 ), true),
						61=> (D_ipd(10)'last_event,  tpd_D_O((511 - 24)- 32*5 ), true),
						62 => (D_ipd(11)'last_event,  tpd_D_O((511 - 24)- 32*4 ), true),
						63 => (D_ipd(12)'last_event,  tpd_D_O((511 - 24)- 32*3 ), true),
						64=> (D_ipd(13)'last_event,  tpd_D_O((511 - 24)- 32*2 ), true),
						65=> (D_ipd(14)'last_event,  tpd_D_O((511 - 24)- 32*1 ), true), 
						66=> (D_ipd(15)'last_event,  tpd_D_O((511 - 24)- 32*0 ), true),
						67=> (CI_ipd'last_event, tpd_CI_O(7), true) ,  
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(7), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(7),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(7),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(7),true)),
      Mode          => VitalTransport,
	  IgnoreDefaultDelay => TRUE,
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);	   
	  
	  
	  	   VitalPathDelay01 (
      OutSignal     => O(8),
      GlitchData    => O_GlitchData(8),
      OutSignalName => "O(8)",
      OutTemp       => O_zd(8),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(8), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(8), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(8), true),
						3 => (A_ipd(0)'last_event,  tpd_A_O((511 - 23)- 32*15 ), true),
						4 => (A_ipd(1)'last_event,  tpd_A_O((511 - 23)- 32*14 ), true),
						5 => (A_ipd(2)'last_event,  tpd_A_O((511 - 23)- 32*13 ), true),
						6 => (A_ipd(3)'last_event,  tpd_A_O((511 - 23)- 32*12 ), true),
						7 => (A_ipd(4)'last_event,  tpd_A_O((511 - 23)- 32*11 ), true), 
						8 => (A_ipd(5)'last_event,  tpd_A_O((511 - 23)- 32*10 ), true),
						9 => (A_ipd(6)'last_event,  tpd_A_O((511 - 23)- 32*9 ), true),
						10 => (A_ipd(7)'last_event,  tpd_A_O((511 - 23)- 32*8 ), true),
						11=> (A_ipd(8)'last_event,  tpd_A_O((511 - 23)- 32*7 ), true),
						12 => (A_ipd(9)'last_event,  tpd_A_O((511 - 23)- 32*6 ), true),
						13 => (A_ipd(10)'last_event,  tpd_A_O((511 - 23)- 32*5 ), true),
						14 => (A_ipd(11)'last_event,  tpd_A_O((511 - 23)- 32*4 ), true),
						15 => (A_ipd(12)'last_event,  tpd_A_O((511 - 23)- 32*3 ), true),
						16=> (A_ipd(13)'last_event,  tpd_A_O((511 - 23)- 32*2), true),
						17=> (A_ipd(14)'last_event,  tpd_A_O((511 - 23)- 32*1 ), true), 
						18=> (A_ipd(15)'last_event,  tpd_A_O((511 - 23)- 32*0 ), true), 
						19=> (B_ipd(0)'last_event,  tpd_B_O((511 - 23)- 32*15 ), true),
						20 => (B_ipd(1)'last_event,  tpd_B_O((511 - 23)- 32*14 ), true),
						21 => (B_ipd(2)'last_event,  tpd_B_O((511 - 23)- 32*13 ), true),
						22 => (B_ipd(3)'last_event,  tpd_B_O((511 - 23)- 32*12 ), true),
						23=> (B_ipd(4)'last_event,  tpd_B_O((511 - 23)- 32*11 ), true), 
						24=> (B_ipd(5)'last_event,  tpd_B_O((511 - 23)- 32*10 ), true),
						25 => (B_ipd(6)'last_event,  tpd_B_O((511 - 23)- 32*9 ), true),
						26 => (B_ipd(7)'last_event,  tpd_B_O((511 - 23)- 32*8 ), true),
						27=> (B_ipd(8)'last_event,  tpd_B_O((511 - 23)- 32*7), true),
						28 => (B_ipd(9)'last_event,  tpd_B_O((511 - 23)- 32*6 ), true),
						29=> (B_ipd(10)'last_event,  tpd_B_O((511 - 23)- 32*5 ), true),
						30 => (B_ipd(11)'last_event,  tpd_B_O((511 - 23)- 32*4 ), true),
						31 => (B_ipd(12)'last_event,  tpd_B_O((511 - 23)- 32*3 ), true),
						32=> (B_ipd(13)'last_event,  tpd_B_O((511 - 23)- 32*2 ), true),
						33=> (B_ipd(14)'last_event,  tpd_B_O((511 - 23)- 32*1 ), true), 
						34=> (B_ipd(15)'last_event,  tpd_B_O((511 - 23)- 32*0 ), true),
						35=> (C_ipd(0)'last_event,  tpd_C_O((511 - 23)- 32*15 ), true),
						36 => (C_ipd(1)'last_event,  tpd_C_O((511 - 23)- 32*14 ), true),
						37 => (C_ipd(2)'last_event,  tpd_C_O((511 - 23)- 32*13 ), true),
						38 => (C_ipd(3)'last_event,  tpd_C_O((511 - 23)- 32*12 ), true),
						39=> (C_ipd(4)'last_event,  tpd_C_O((511 - 23)- 32*11 ), true), 
						40=> (C_ipd(5)'last_event,  tpd_C_O((511 - 23)- 32*10 ), true),
						41 => (C_ipd(6)'last_event,  tpd_C_O((511 - 23)- 32*9 ), true),
						42 => (C_ipd(7)'last_event,  tpd_C_O((511 - 23)- 32*8 ), true),
						43=> (C_ipd(8)'last_event,  tpd_C_O((511 - 23)- 32*7), true),
						44 => (C_ipd(9)'last_event,  tpd_C_O((511 - 23)- 32*6 ), true),
						45=> (C_ipd(10)'last_event,  tpd_C_O((511 - 23)- 32*5 ), true),
						46 => (C_ipd(11)'last_event,  tpd_C_O((511 - 23)- 32*4 ), true),
						47 => (C_ipd(12)'last_event,  tpd_C_O((511 - 23)- 32*3 ), true),
						48=> (C_ipd(13)'last_event,  tpd_C_O((511 - 23)- 32*2 ), true),
						49=> (C_ipd(14)'last_event,  tpd_C_O((511 - 23)- 32*1 ), true), 
						50=> (C_ipd(15)'last_event,  tpd_C_O((511 - 23)- 32*0 ), true),
						51=> (D_ipd(0)'last_event,  tpd_D_O((511 - 23)- 32*15 ), true),
						52 => (D_ipd(1)'last_event,  tpd_D_O((511 - 23)- 32*14 ), true),
						53 => (D_ipd(2)'last_event,  tpd_D_O((511 - 23)- 32*13 ), true),
						54 => (D_ipd(3)'last_event,  tpd_D_O((511 - 23)- 32*12 ), true),
						55=> (D_ipd(4)'last_event,  tpd_D_O((511 - 23)- 32*11 ), true), 
						56=> (D_ipd(5)'last_event,  tpd_D_O((511 - 23)- 32*10 ), true),
						57 => (D_ipd(6)'last_event,  tpd_D_O((511 - 23)- 32*9 ), true),
						58 => (D_ipd(7)'last_event,  tpd_D_O((511 - 23)- 32*8 ), true),
						59=> (D_ipd(8)'last_event,  tpd_D_O((511 - 23)- 32*7 ), true),
						60 => (D_ipd(9)'last_event,  tpd_D_O((511 - 23)- 32*6 ), true),
						61=> (D_ipd(10)'last_event,  tpd_D_O((511 - 23)- 32*5 ), true),
						62 => (D_ipd(11)'last_event,  tpd_D_O((511 - 23)- 32*4 ), true),
						63 => (D_ipd(12)'last_event,  tpd_D_O((511 - 23)- 32*3 ), true),
						64=> (D_ipd(13)'last_event,  tpd_D_O((511 - 23)- 32*2 ), true),
						65=> (D_ipd(14)'last_event,  tpd_D_O((511 - 23)- 32*1 ), true), 
						66=> (D_ipd(15)'last_event,  tpd_D_O((511 - 23)- 32*0 ), true),
						67=> (CI_ipd'last_event, tpd_CI_O(8), true)  ,  
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(8), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(8),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(8),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(8),true)),
      Mode          => VitalTransport,	
	  IgnoreDefaultDelay => TRUE, 
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);
	  
	  
	  	   VitalPathDelay01 (
      OutSignal     => O(9),
      GlitchData    => O_GlitchData(9),
      OutSignalName => "O(9)",
      OutTemp       => O_zd(9),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(9), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(9), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(9), true),
							3 => (A_ipd(0)'last_event,  tpd_A_O((511 - 22)- 32*15 ), true),
						4 => (A_ipd(1)'last_event,  tpd_A_O((511 - 22)- 32*14 ), true),
						5 => (A_ipd(2)'last_event,  tpd_A_O((511 - 22)- 32*13 ), true),
						6 => (A_ipd(3)'last_event,  tpd_A_O((511 - 22)- 32*12 ), true),
						7 => (A_ipd(4)'last_event,  tpd_A_O((511 - 22)- 32*11 ), true), 
						8 => (A_ipd(5)'last_event,  tpd_A_O((511 - 22)- 32*10 ), true),
						9 => (A_ipd(6)'last_event,  tpd_A_O((511 - 22)- 32*9 ), true),
						10 => (A_ipd(7)'last_event,  tpd_A_O((511 - 22)- 32*8 ), true),
						11=> (A_ipd(8)'last_event,  tpd_A_O((511 - 22)- 32*7 ), true),
						12 => (A_ipd(9)'last_event,  tpd_A_O((511 - 22)- 32*6 ), true),
						13 => (A_ipd(10)'last_event,  tpd_A_O((511 - 22)- 32*5 ), true),
						14 => (A_ipd(11)'last_event,  tpd_A_O((511 - 22)- 32*4 ), true),
						15 => (A_ipd(12)'last_event,  tpd_A_O((511 - 22)- 32*3 ), true),
						16=> (A_ipd(13)'last_event,  tpd_A_O((511 - 22)- 32*2), true),
						17=> (A_ipd(14)'last_event,  tpd_A_O((511 - 22)- 32*1 ), true), 
						18=> (A_ipd(15)'last_event,  tpd_A_O((511 - 22)- 32*0 ), true), 
						19=> (B_ipd(0)'last_event,  tpd_B_O((511 - 22)- 32*15 ), true),
						20 => (B_ipd(1)'last_event,  tpd_B_O((511 - 22)- 32*14 ), true),
						21 => (B_ipd(2)'last_event,  tpd_B_O((511 - 22)- 32*13 ), true),
						22 => (B_ipd(3)'last_event,  tpd_B_O((511 - 22)- 32*12 ), true),
						23=> (B_ipd(4)'last_event,  tpd_B_O((511 - 22)- 32*11 ), true), 
						24=> (B_ipd(5)'last_event,  tpd_B_O((511 - 22)- 32*10 ), true),
						25 => (B_ipd(6)'last_event,  tpd_B_O((511 - 22)- 32*9 ), true),
						26 => (B_ipd(7)'last_event,  tpd_B_O((511 - 22)- 32*8 ), true),
						27=> (B_ipd(8)'last_event,  tpd_B_O((511 - 22)- 32*7), true),
						28 => (B_ipd(9)'last_event,  tpd_B_O((511 - 22)- 32*6 ), true),
						29=> (B_ipd(10)'last_event,  tpd_B_O((511 - 22)- 32*5 ), true),
						30 => (B_ipd(11)'last_event,  tpd_B_O((511 - 22)- 32*4 ), true),
						31 => (B_ipd(12)'last_event,  tpd_B_O((511 - 22)- 32*3 ), true),
						32=> (B_ipd(13)'last_event,  tpd_B_O((511 - 22)- 32*2 ), true),
						33=> (B_ipd(14)'last_event,  tpd_B_O((511 - 22)- 32*1 ), true), 
						34=> (B_ipd(15)'last_event,  tpd_B_O((511 - 22)- 32*0 ), true),
						35=> (C_ipd(0)'last_event,  tpd_C_O((511 - 22)- 32*15 ), true),
						36 => (C_ipd(1)'last_event,  tpd_C_O((511 - 22)- 32*14 ), true),
						37 => (C_ipd(2)'last_event,  tpd_C_O((511 - 22)- 32*13 ), true),
						38 => (C_ipd(3)'last_event,  tpd_C_O((511 - 22)- 32*12 ), true),
						39=> (C_ipd(4)'last_event,  tpd_C_O((511 - 22)- 32*11 ), true), 
						40=> (C_ipd(5)'last_event,  tpd_C_O((511 - 22)- 32*10 ), true),
						41 => (C_ipd(6)'last_event,  tpd_C_O((511 - 22)- 32*9 ), true),
						42 => (C_ipd(7)'last_event,  tpd_C_O((511 - 22)- 32*8 ), true),
						43=> (C_ipd(8)'last_event,  tpd_C_O((511 - 22)- 32*7), true),
						44 => (C_ipd(9)'last_event,  tpd_C_O((511 - 22)- 32*6 ), true),
						45=> (C_ipd(10)'last_event,  tpd_C_O((511 - 22)- 32*5 ), true),
						46 => (C_ipd(11)'last_event,  tpd_C_O((511 - 22)- 32*4 ), true),
						47 => (C_ipd(12)'last_event,  tpd_C_O((511 - 22)- 32*3 ), true),
						48=> (C_ipd(13)'last_event,  tpd_C_O((511 - 22)- 32*2 ), true),
						49=> (C_ipd(14)'last_event,  tpd_C_O((511 - 22)- 32*1 ), true), 
						50=> (C_ipd(15)'last_event,  tpd_C_O((511 - 22)- 32*0 ), true),
						51=> (D_ipd(0)'last_event,  tpd_D_O((511 - 22)- 32*15 ), true),
						52 => (D_ipd(1)'last_event,  tpd_D_O((511 - 22)- 32*14 ), true),
						53 => (D_ipd(2)'last_event,  tpd_D_O((511 - 22)- 32*13 ), true),
						54 => (D_ipd(3)'last_event,  tpd_D_O((511 - 22)- 32*12 ), true),
						55=> (D_ipd(4)'last_event,  tpd_D_O((511 - 22)- 32*11 ), true), 
						56=> (D_ipd(5)'last_event,  tpd_D_O((511 - 22)- 32*10 ), true),
						57 => (D_ipd(6)'last_event,  tpd_D_O((511 - 22)- 32*9 ), true),
						58 => (D_ipd(7)'last_event,  tpd_D_O((511 - 22)- 32*8 ), true),
						59=> (D_ipd(8)'last_event,  tpd_D_O((511 - 22)- 32*7 ), true),
						60 => (D_ipd(9)'last_event,  tpd_D_O((511 - 22)- 32*6 ), true),
						61=> (D_ipd(10)'last_event,  tpd_D_O((511 - 22)- 32*5 ), true),
						62 => (D_ipd(11)'last_event,  tpd_D_O((511 - 22)- 32*4 ), true),
						63 => (D_ipd(12)'last_event,  tpd_D_O((511 - 22)- 32*3 ), true),
						64=> (D_ipd(13)'last_event,  tpd_D_O((511 - 22)- 32*2 ), true),
						65=> (D_ipd(14)'last_event,  tpd_D_O((511 - 22)- 32*1 ), true), 
						66=> (D_ipd(15)'last_event,  tpd_D_O((511 - 22)- 32*0 ), true),
						67=> (CI_ipd'last_event, tpd_CI_O(9), true)  ,  
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(9), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(9),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(9),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(9),true)),
      Mode          => VitalTransport, 
	  IgnoreDefaultDelay => TRUE,
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);
	  
	  
	  	   VitalPathDelay01 (
      OutSignal     => O(10),
      GlitchData    => O_GlitchData(10),
      OutSignalName => "O(10)",
      OutTemp       => O_zd(10),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(10), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(10), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(10), true),
							3 => (A_ipd(0)'last_event,  tpd_A_O((511 - 21)- 32*15 ), true),
						4 => (A_ipd(1)'last_event,  tpd_A_O((511 - 21)- 32*14 ), true),
						5 => (A_ipd(2)'last_event,  tpd_A_O((511 - 21)- 32*13 ), true),
						6 => (A_ipd(3)'last_event,  tpd_A_O((511 - 21)- 32*12 ), true),
						7 => (A_ipd(4)'last_event,  tpd_A_O((511 - 21)- 32*11 ), true), 
						8 => (A_ipd(5)'last_event,  tpd_A_O((511 - 21)- 32*10 ), true),
						9 => (A_ipd(6)'last_event,  tpd_A_O((511 - 21)- 32*9 ), true),
						10 => (A_ipd(7)'last_event,  tpd_A_O((511 - 21)- 32*8 ), true),
						11=> (A_ipd(8)'last_event,  tpd_A_O((511 - 21)- 32*7 ), true),
						12 => (A_ipd(9)'last_event,  tpd_A_O((511 - 21)- 32*6 ), true),
						13 => (A_ipd(10)'last_event,  tpd_A_O((511 - 21)- 32*5 ), true),
						14 => (A_ipd(11)'last_event,  tpd_A_O((511 - 21)- 32*4 ), true),
						15 => (A_ipd(12)'last_event,  tpd_A_O((511 - 21)- 32*3 ), true),
						16=> (A_ipd(13)'last_event,  tpd_A_O((511 - 21)- 32*2), true),
						17=> (A_ipd(14)'last_event,  tpd_A_O((511 - 21)- 32*1 ), true), 
						18=> (A_ipd(15)'last_event,  tpd_A_O((511 - 21)- 32*0 ), true), 
						19=> (B_ipd(0)'last_event,  tpd_B_O((511 - 21)- 32*15 ), true),
						20 => (B_ipd(1)'last_event,  tpd_B_O((511 - 21)- 32*14 ), true),
						21 => (B_ipd(2)'last_event,  tpd_B_O((511 - 21)- 32*13 ), true),
						22 => (B_ipd(3)'last_event,  tpd_B_O((511 - 21)- 32*12 ), true),
						23=> (B_ipd(4)'last_event,  tpd_B_O((511 - 21)- 32*11 ), true), 
						24=> (B_ipd(5)'last_event,  tpd_B_O((511 - 21)- 32*10 ), true),
						25 => (B_ipd(6)'last_event,  tpd_B_O((511 - 21)- 32*9 ), true),
						26 => (B_ipd(7)'last_event,  tpd_B_O((511 - 21)- 32*8 ), true),
						27=> (B_ipd(8)'last_event,  tpd_B_O((511 - 21)- 32*7), true),
						28 => (B_ipd(9)'last_event,  tpd_B_O((511 - 21)- 32*6 ), true),
						29=> (B_ipd(10)'last_event,  tpd_B_O((511 - 21)- 32*5 ), true),
						30 => (B_ipd(11)'last_event,  tpd_B_O((511 - 21)- 32*4 ), true),
						31 => (B_ipd(12)'last_event,  tpd_B_O((511 - 21)- 32*3 ), true),
						32=> (B_ipd(13)'last_event,  tpd_B_O((511 - 21)- 32*2 ), true),
						33=> (B_ipd(14)'last_event,  tpd_B_O((511 - 21)- 32*1 ), true), 
						34=> (B_ipd(15)'last_event,  tpd_B_O((511 - 21)- 32*0 ), true),
						35=> (C_ipd(0)'last_event,  tpd_C_O((511 - 21)- 32*15 ), true),
						36 => (C_ipd(1)'last_event,  tpd_C_O((511 - 21)- 32*14 ), true),
						37 => (C_ipd(2)'last_event,  tpd_C_O((511 - 21)- 32*13 ), true),
						38 => (C_ipd(3)'last_event,  tpd_C_O((511 - 21)- 32*12 ), true),
						39=> (C_ipd(4)'last_event,  tpd_C_O((511 - 21)- 32*11 ), true), 
						40=> (C_ipd(5)'last_event,  tpd_C_O((511 - 21)- 32*10 ), true),
						41 => (C_ipd(6)'last_event,  tpd_C_O((511 - 21)- 32*9 ), true),
						42 => (C_ipd(7)'last_event,  tpd_C_O((511 - 21)- 32*8 ), true),
						43=> (C_ipd(8)'last_event,  tpd_C_O((511 - 21)- 32*7), true),
						44 => (C_ipd(9)'last_event,  tpd_C_O((511 - 21)- 32*6 ), true),
						45=> (C_ipd(10)'last_event,  tpd_C_O((511 - 21)- 32*5 ), true),
						46 => (C_ipd(11)'last_event,  tpd_C_O((511 - 21)- 32*4 ), true),
						47 => (C_ipd(12)'last_event,  tpd_C_O((511 - 21)- 32*3 ), true),
						48=> (C_ipd(13)'last_event,  tpd_C_O((511 - 21)- 32*2 ), true),
						49=> (C_ipd(14)'last_event,  tpd_C_O((511 - 21)- 32*1 ), true), 
						50=> (C_ipd(15)'last_event,  tpd_C_O((511 - 21)- 32*0 ), true),
						51=> (D_ipd(0)'last_event,  tpd_D_O((511 - 21)- 32*15 ), true),
						52 => (D_ipd(1)'last_event,  tpd_D_O((511 - 21)- 32*14 ), true),
						53 => (D_ipd(2)'last_event,  tpd_D_O((511 - 21)- 32*13 ), true),
						54 => (D_ipd(3)'last_event,  tpd_D_O((511 - 21)- 32*12 ), true),
						55=> (D_ipd(4)'last_event,  tpd_D_O((511 - 21)- 32*11 ), true), 
						56=> (D_ipd(5)'last_event,  tpd_D_O((511 - 21)- 32*10 ), true),
						57 => (D_ipd(6)'last_event,  tpd_D_O((511 - 21)- 32*9 ), true),
						58 => (D_ipd(7)'last_event,  tpd_D_O((511 - 21)- 32*8 ), true),
						59=> (D_ipd(8)'last_event,  tpd_D_O((511 - 21)- 32*7 ), true),
						60 => (D_ipd(9)'last_event,  tpd_D_O((511 - 21)- 32*6 ), true),
						61=> (D_ipd(10)'last_event,  tpd_D_O((511 - 21)- 32*5 ), true),
						62 => (D_ipd(11)'last_event,  tpd_D_O((511 - 21)- 32*4 ), true),
						63 => (D_ipd(12)'last_event,  tpd_D_O((511 - 21)- 32*3 ), true),
						64=> (D_ipd(13)'last_event,  tpd_D_O((511 - 21)- 32*2 ), true),
						65=> (D_ipd(14)'last_event,  tpd_D_O((511 - 21)- 32*1 ), true), 
						66=> (D_ipd(15)'last_event,  tpd_D_O((511 - 21)- 32*0 ), true),
						67=> (CI_ipd'last_event, tpd_CI_O(10), true) ,  
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(10), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(10),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(10),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(10),true)),
      Mode          => VitalTransport,
	  IgnoreDefaultDelay => TRUE, 
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);
	  
	
	
	  	   VitalPathDelay01 (
      OutSignal     => O(11),
      GlitchData    => O_GlitchData(11),
      OutSignalName => "O(11)",
      OutTemp       => O_zd(11),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(11), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(11), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(11), true),
							3 => (A_ipd(0)'last_event,  tpd_A_O((511 - 20)- 32*15 ), true),
						4 => (A_ipd(1)'last_event,  tpd_A_O((511 - 20)- 32*14 ), true),
						5 => (A_ipd(2)'last_event,  tpd_A_O((511 - 20)- 32*13 ), true),
						6 => (A_ipd(3)'last_event,  tpd_A_O((511 - 20)- 32*12 ), true),
						7 => (A_ipd(4)'last_event,  tpd_A_O((511 - 20)- 32*11 ), true), 
						8 => (A_ipd(5)'last_event,  tpd_A_O((511 - 20)- 32*10 ), true),
						9 => (A_ipd(6)'last_event,  tpd_A_O((511 - 20)- 32*9 ), true),
						10 => (A_ipd(7)'last_event,  tpd_A_O((511 - 20)- 32*8 ), true),
						11=> (A_ipd(8)'last_event,  tpd_A_O((511 - 20)- 32*7 ), true),
						12 => (A_ipd(9)'last_event,  tpd_A_O((511 - 20)- 32*6 ), true),
						13 => (A_ipd(10)'last_event,  tpd_A_O((511 - 20)- 32*5 ), true),
						14 => (A_ipd(11)'last_event,  tpd_A_O((511 - 20)- 32*4 ), true),
						15 => (A_ipd(12)'last_event,  tpd_A_O((511 - 20)- 32*3 ), true),
						16=> (A_ipd(13)'last_event,  tpd_A_O((511 - 20)- 32*2), true),
						17=> (A_ipd(14)'last_event,  tpd_A_O((511 - 20)- 32*1 ), true), 
						18=> (A_ipd(15)'last_event,  tpd_A_O((511 - 20)- 32*0 ), true), 
						19=> (B_ipd(0)'last_event,  tpd_B_O((511 - 20)- 32*15 ), true),
						20 => (B_ipd(1)'last_event,  tpd_B_O((511 - 20)- 32*14 ), true),
						21 => (B_ipd(2)'last_event,  tpd_B_O((511 - 20)- 32*13 ), true),
						22 => (B_ipd(3)'last_event,  tpd_B_O((511 - 20)- 32*12 ), true),
						23=> (B_ipd(4)'last_event,  tpd_B_O((511 - 20)- 32*11 ), true), 
						24=> (B_ipd(5)'last_event,  tpd_B_O((511 - 20)- 32*10 ), true),
						25 => (B_ipd(6)'last_event,  tpd_B_O((511 - 20)- 32*9 ), true),
						26 => (B_ipd(7)'last_event,  tpd_B_O((511 - 20)- 32*8 ), true),
						27=> (B_ipd(8)'last_event,  tpd_B_O((511 - 20)- 32*7), true),
						28 => (B_ipd(9)'last_event,  tpd_B_O((511 - 20)- 32*6 ), true),
						29=> (B_ipd(10)'last_event,  tpd_B_O((511 - 20)- 32*5 ), true),
						30 => (B_ipd(11)'last_event,  tpd_B_O((511 - 20)- 32*4 ), true),
						31 => (B_ipd(12)'last_event,  tpd_B_O((511 - 20)- 32*3 ), true),
						32=> (B_ipd(13)'last_event,  tpd_B_O((511 - 20)- 32*2 ), true),
						33=> (B_ipd(14)'last_event,  tpd_B_O((511 - 20)- 32*1 ), true), 
						34=> (B_ipd(15)'last_event,  tpd_B_O((511 - 20)- 32*0 ), true),
						35=> (C_ipd(0)'last_event,  tpd_C_O((511 - 20)- 32*15 ), true),
						36 => (C_ipd(1)'last_event,  tpd_C_O((511 - 20)- 32*14 ), true),
						37 => (C_ipd(2)'last_event,  tpd_C_O((511 - 20)- 32*13 ), true),
						38 => (C_ipd(3)'last_event,  tpd_C_O((511 - 20)- 32*12 ), true),
						39=> (C_ipd(4)'last_event,  tpd_C_O((511 - 20)- 32*11 ), true), 
						40=> (C_ipd(5)'last_event,  tpd_C_O((511 - 20)- 32*10 ), true),
						41 => (C_ipd(6)'last_event,  tpd_C_O((511 - 20)- 32*9 ), true),
						42 => (C_ipd(7)'last_event,  tpd_C_O((511 - 20)- 32*8 ), true),
						43=> (C_ipd(8)'last_event,  tpd_C_O((511 - 20)- 32*7), true),
						44 => (C_ipd(9)'last_event,  tpd_C_O((511 - 20)- 32*6 ), true),
						45=> (C_ipd(10)'last_event,  tpd_C_O((511 - 20)- 32*5 ), true),
						46 => (C_ipd(11)'last_event,  tpd_C_O((511 - 20)- 32*4 ), true),
						47 => (C_ipd(12)'last_event,  tpd_C_O((511 - 20)- 32*3 ), true),
						48=> (C_ipd(13)'last_event,  tpd_C_O((511 - 20)- 32*2 ), true),
						49=> (C_ipd(14)'last_event,  tpd_C_O((511 - 20)- 32*1 ), true), 
						50=> (C_ipd(15)'last_event,  tpd_C_O((511 - 20)- 32*0 ), true),
						51=> (D_ipd(0)'last_event,  tpd_D_O((511 - 20)- 32*15 ), true),
						52 => (D_ipd(1)'last_event,  tpd_D_O((511 - 20)- 32*14 ), true),
						53 => (D_ipd(2)'last_event,  tpd_D_O((511 - 20)- 32*13 ), true),
						54 => (D_ipd(3)'last_event,  tpd_D_O((511 - 20)- 32*12 ), true),
						55=> (D_ipd(4)'last_event,  tpd_D_O((511 - 20)- 32*11 ), true), 
						56=> (D_ipd(5)'last_event,  tpd_D_O((511 - 20)- 32*10 ), true),
						57 => (D_ipd(6)'last_event,  tpd_D_O((511 - 20)- 32*9 ), true),
						58 => (D_ipd(7)'last_event,  tpd_D_O((511 - 20)- 32*8 ), true),
						59=> (D_ipd(8)'last_event,  tpd_D_O((511 - 20)- 32*7 ), true),
						60 => (D_ipd(9)'last_event,  tpd_D_O((511 - 20)- 32*6 ), true),
						61=> (D_ipd(10)'last_event,  tpd_D_O((511 - 20)- 32*5 ), true),
						62 => (D_ipd(11)'last_event,  tpd_D_O((511 - 20)- 32*4 ), true),
						63 => (D_ipd(12)'last_event,  tpd_D_O((511 - 20)- 32*3 ), true),
						64=> (D_ipd(13)'last_event,  tpd_D_O((511 - 20)- 32*2 ), true),
						65=> (D_ipd(14)'last_event,  tpd_D_O((511 - 20)- 32*1 ), true), 
						66=> (D_ipd(15)'last_event,  tpd_D_O((511 - 20)- 32*0 ), true),
						67=> (CI_ipd'last_event, tpd_CI_O(11), true)  ,  
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(11), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(11),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(11),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(11),true)),
      Mode          => VitalTransport,		  
	  IgnoreDefaultDelay => TRUE, 
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);	 
	  
	  
	  	   VitalPathDelay01 (
      OutSignal     => O(12),
      GlitchData    => O_GlitchData(12),
      OutSignalName => "O(12)",
      OutTemp       => O_zd(12),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(12), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(12), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(12), true),
							3 => (A_ipd(0)'last_event,  tpd_A_O((511 - 19)- 32*15 ), true),
						4 => (A_ipd(1)'last_event,  tpd_A_O((511 - 19)- 32*14 ), true),
						5 => (A_ipd(2)'last_event,  tpd_A_O((511 - 19)- 32*13 ), true),
						6 => (A_ipd(3)'last_event,  tpd_A_O((511 - 19)- 32*12 ), true),
						7 => (A_ipd(4)'last_event,  tpd_A_O((511 - 19)- 32*11 ), true), 
						8 => (A_ipd(5)'last_event,  tpd_A_O((511 - 19)- 32*10 ), true),
						9 => (A_ipd(6)'last_event,  tpd_A_O((511 - 19)- 32*9 ), true),
						10 => (A_ipd(7)'last_event,  tpd_A_O((511 - 19)- 32*8 ), true),
						11=> (A_ipd(8)'last_event,  tpd_A_O((511 - 19)- 32*7 ), true),
						12 => (A_ipd(9)'last_event,  tpd_A_O((511 - 19)- 32*6 ), true),
						13 => (A_ipd(10)'last_event,  tpd_A_O((511 - 19)- 32*5 ), true),
						14 => (A_ipd(11)'last_event,  tpd_A_O((511 - 19)- 32*4 ), true),
						15 => (A_ipd(12)'last_event,  tpd_A_O((511 - 19)- 32*3 ), true),
						16=> (A_ipd(13)'last_event,  tpd_A_O((511 - 19)- 32*2), true),
						17=> (A_ipd(14)'last_event,  tpd_A_O((511 - 19)- 32*1 ), true), 
						18=> (A_ipd(15)'last_event,  tpd_A_O((511 - 19)- 32*0 ), true), 
						19=> (B_ipd(0)'last_event,  tpd_B_O((511 - 19)- 32*15 ), true),
						20 => (B_ipd(1)'last_event,  tpd_B_O((511 - 19)- 32*14 ), true),
						21 => (B_ipd(2)'last_event,  tpd_B_O((511 - 19)- 32*13 ), true),
						22 => (B_ipd(3)'last_event,  tpd_B_O((511 - 19)- 32*12 ), true),
						23=> (B_ipd(4)'last_event,  tpd_B_O((511 - 19)- 32*11 ), true), 
						24=> (B_ipd(5)'last_event,  tpd_B_O((511 - 19)- 32*10 ), true),
						25 => (B_ipd(6)'last_event,  tpd_B_O((511 - 19)- 32*9 ), true),
						26 => (B_ipd(7)'last_event,  tpd_B_O((511 - 19)- 32*8 ), true),
						27=> (B_ipd(8)'last_event,  tpd_B_O((511 - 19)- 32*7), true),
						28 => (B_ipd(9)'last_event,  tpd_B_O((511 - 19)- 32*6 ), true),
						29=> (B_ipd(10)'last_event,  tpd_B_O((511 - 19)- 32*5 ), true),
						30 => (B_ipd(11)'last_event,  tpd_B_O((511 - 19)- 32*4 ), true),
						31 => (B_ipd(12)'last_event,  tpd_B_O((511 - 19)- 32*3 ), true),
						32=> (B_ipd(13)'last_event,  tpd_B_O((511 - 19)- 32*2 ), true),
						33=> (B_ipd(14)'last_event,  tpd_B_O((511 - 19)- 32*1 ), true), 
						34=> (B_ipd(15)'last_event,  tpd_B_O((511 - 19)- 32*0 ), true),
						35=> (C_ipd(0)'last_event,  tpd_C_O((511 - 19)- 32*15 ), true),
						36 => (C_ipd(1)'last_event,  tpd_C_O((511 - 19)- 32*14 ), true),
						37 => (C_ipd(2)'last_event,  tpd_C_O((511 - 19)- 32*13 ), true),
						38 => (C_ipd(3)'last_event,  tpd_C_O((511 - 19)- 32*12 ), true),
						39=> (C_ipd(4)'last_event,  tpd_C_O((511 - 19)- 32*11 ), true), 
						40=> (C_ipd(5)'last_event,  tpd_C_O((511 - 19)- 32*10 ), true),
						41 => (C_ipd(6)'last_event,  tpd_C_O((511 - 19)- 32*9 ), true),
						42 => (C_ipd(7)'last_event,  tpd_C_O((511 - 19)- 32*8 ), true),
						43=> (C_ipd(8)'last_event,  tpd_C_O((511 - 19)- 32*7), true),
						44 => (C_ipd(9)'last_event,  tpd_C_O((511 - 19)- 32*6 ), true),
						45=> (C_ipd(10)'last_event,  tpd_C_O((511 - 19)- 32*5 ), true),
						46 => (C_ipd(11)'last_event,  tpd_C_O((511 - 19)- 32*4 ), true),
						47 => (C_ipd(12)'last_event,  tpd_C_O((511 - 19)- 32*3 ), true),
						48=> (C_ipd(13)'last_event,  tpd_C_O((511 - 19)- 32*2 ), true),
						49=> (C_ipd(14)'last_event,  tpd_C_O((511 - 19)- 32*1 ), true), 
						50=> (C_ipd(15)'last_event,  tpd_C_O((511 - 19)- 32*0 ), true),
						51=> (D_ipd(0)'last_event,  tpd_D_O((511 - 19)- 32*15 ), true),
						52 => (D_ipd(1)'last_event,  tpd_D_O((511 - 19)- 32*14 ), true),
						53 => (D_ipd(2)'last_event,  tpd_D_O((511 - 19)- 32*13 ), true),
						54 => (D_ipd(3)'last_event,  tpd_D_O((511 - 19)- 32*12 ), true),
						55=> (D_ipd(4)'last_event,  tpd_D_O((511 - 19)- 32*11 ), true), 
						56=> (D_ipd(5)'last_event,  tpd_D_O((511 - 19)- 32*10 ), true),
						57 => (D_ipd(6)'last_event,  tpd_D_O((511 - 19)- 32*9 ), true),
						58 => (D_ipd(7)'last_event,  tpd_D_O((511 - 19)- 32*8 ), true),
						59=> (D_ipd(8)'last_event,  tpd_D_O((511 - 19)- 32*7 ), true),
						60 => (D_ipd(9)'last_event,  tpd_D_O((511 - 19)- 32*6 ), true),
						61=> (D_ipd(10)'last_event,  tpd_D_O((511 - 19)- 32*5 ), true),
						62 => (D_ipd(11)'last_event,  tpd_D_O((511 - 19)- 32*4 ), true),
						63 => (D_ipd(12)'last_event,  tpd_D_O((511 - 19)- 32*3 ), true),
						64=> (D_ipd(13)'last_event,  tpd_D_O((511 - 19)- 32*2 ), true),
						65=> (D_ipd(14)'last_event,  tpd_D_O((511 - 19)- 32*1 ), true), 
						66=> (D_ipd(15)'last_event,  tpd_D_O((511 - 19)- 32*0 ), true),
						67=> (CI_ipd'last_event, tpd_CI_O(12), true)  ,  
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(12), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(12),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(12),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(12),true)),
      Mode          => VitalTransport, 
	  IgnoreDefaultDelay => TRUE,
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);				   
	  
	  
	  	   VitalPathDelay01 (
      OutSignal     => O(13),
      GlitchData    => O_GlitchData(13),
      OutSignalName => "O(13)",
      OutTemp       => O_zd(13),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(13), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(13), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(13), true),
						3 => (A_ipd(0)'last_event,  tpd_A_O((511 - 18)- 32*15 ), true),
						4 => (A_ipd(1)'last_event,  tpd_A_O((511 - 18)- 32*14 ), true),
						5 => (A_ipd(2)'last_event,  tpd_A_O((511 - 18)- 32*13 ), true),
						6 => (A_ipd(3)'last_event,  tpd_A_O((511 - 18)- 32*12 ), true),
						7 => (A_ipd(4)'last_event,  tpd_A_O((511 - 18)- 32*11 ), true), 
						8 => (A_ipd(5)'last_event,  tpd_A_O((511 - 18)- 32*10 ), true),
						9 => (A_ipd(6)'last_event,  tpd_A_O((511 - 18)- 32*9 ), true),
						10 => (A_ipd(7)'last_event,  tpd_A_O((511 - 18)- 32*8 ), true),
						11=> (A_ipd(8)'last_event,  tpd_A_O((511 - 18)- 32*7 ), true),
						12 => (A_ipd(9)'last_event,  tpd_A_O((511 - 18)- 32*6 ), true),
						13 => (A_ipd(10)'last_event,  tpd_A_O((511 - 18)- 32*5 ), true),
						14 => (A_ipd(11)'last_event,  tpd_A_O((511 - 18)- 32*4 ), true),
						15 => (A_ipd(12)'last_event,  tpd_A_O((511 - 18)- 32*3 ), true),
						16=> (A_ipd(13)'last_event,  tpd_A_O((511 - 18)- 32*2), true),
						17=> (A_ipd(14)'last_event,  tpd_A_O((511 - 18)- 32*1 ), true), 
						18=> (A_ipd(15)'last_event,  tpd_A_O((511 - 18)- 32*0 ), true), 
						19=> (B_ipd(0)'last_event,  tpd_B_O((511 - 18)- 32*15 ), true),
						20 => (B_ipd(1)'last_event,  tpd_B_O((511 - 18)- 32*14 ), true),
						21 => (B_ipd(2)'last_event,  tpd_B_O((511 - 18)- 32*13 ), true),
						22 => (B_ipd(3)'last_event,  tpd_B_O((511 - 18)- 32*12 ), true),
						23=> (B_ipd(4)'last_event,  tpd_B_O((511 - 18)- 32*11 ), true), 
						24=> (B_ipd(5)'last_event,  tpd_B_O((511 - 18)- 32*10 ), true),
						25 => (B_ipd(6)'last_event,  tpd_B_O((511 - 18)- 32*9 ), true),
						26 => (B_ipd(7)'last_event,  tpd_B_O((511 - 18)- 32*8 ), true),
						27=> (B_ipd(8)'last_event,  tpd_B_O((511 - 18)- 32*7), true),
						28 => (B_ipd(9)'last_event,  tpd_B_O((511 - 18)- 32*6 ), true),
						29=> (B_ipd(10)'last_event,  tpd_B_O((511 - 18)- 32*5 ), true),
						30 => (B_ipd(11)'last_event,  tpd_B_O((511 - 18)- 32*4 ), true),
						31 => (B_ipd(12)'last_event,  tpd_B_O((511 - 18)- 32*3 ), true),
						32=> (B_ipd(13)'last_event,  tpd_B_O((511 - 18)- 32*2 ), true),
						33=> (B_ipd(14)'last_event,  tpd_B_O((511 - 18)- 32*1 ), true), 
						34=> (B_ipd(15)'last_event,  tpd_B_O((511 - 18)- 32*0 ), true),
						35=> (C_ipd(0)'last_event,  tpd_C_O((511 - 18)- 32*15 ), true),
						36 => (C_ipd(1)'last_event,  tpd_C_O((511 - 18)- 32*14 ), true),
						37 => (C_ipd(2)'last_event,  tpd_C_O((511 - 18)- 32*13 ), true),
						38 => (C_ipd(3)'last_event,  tpd_C_O((511 - 18)- 32*12 ), true),
						39=> (C_ipd(4)'last_event,  tpd_C_O((511 - 18)- 32*11 ), true), 
						40=> (C_ipd(5)'last_event,  tpd_C_O((511 - 18)- 32*10 ), true),
						41 => (C_ipd(6)'last_event,  tpd_C_O((511 - 18)- 32*9 ), true),
						42 => (C_ipd(7)'last_event,  tpd_C_O((511 - 18)- 32*8 ), true),
						43=> (C_ipd(8)'last_event,  tpd_C_O((511 - 18)- 32*7), true),
						44 => (C_ipd(9)'last_event,  tpd_C_O((511 - 18)- 32*6 ), true),
						45=> (C_ipd(10)'last_event,  tpd_C_O((511 - 18)- 32*5 ), true),
						46 => (C_ipd(11)'last_event,  tpd_C_O((511 - 18)- 32*4 ), true),
						47 => (C_ipd(12)'last_event,  tpd_C_O((511 - 18)- 32*3 ), true),
						48=> (C_ipd(13)'last_event,  tpd_C_O((511 - 18)- 32*2 ), true),
						49=> (C_ipd(14)'last_event,  tpd_C_O((511 - 18)- 32*1 ), true), 
						50=> (C_ipd(15)'last_event,  tpd_C_O((511 - 18)- 32*0 ), true),
						51=> (D_ipd(0)'last_event,  tpd_D_O((511 - 18)- 32*15 ), true),
						52 => (D_ipd(1)'last_event,  tpd_D_O((511 - 18)- 32*14 ), true),
						53 => (D_ipd(2)'last_event,  tpd_D_O((511 - 18)- 32*13 ), true),
						54 => (D_ipd(3)'last_event,  tpd_D_O((511 - 18)- 32*12 ), true),
						55=> (D_ipd(4)'last_event,  tpd_D_O((511 - 18)- 32*11 ), true), 
						56=> (D_ipd(5)'last_event,  tpd_D_O((511 - 18)- 32*10 ), true),
						57 => (D_ipd(6)'last_event,  tpd_D_O((511 - 18)- 32*9 ), true),
						58 => (D_ipd(7)'last_event,  tpd_D_O((511 - 18)- 32*8 ), true),
						59=> (D_ipd(8)'last_event,  tpd_D_O((511 - 18)- 32*7 ), true),
						60 => (D_ipd(9)'last_event,  tpd_D_O((511 - 18)- 32*6 ), true),
						61=> (D_ipd(10)'last_event,  tpd_D_O((511 - 18)- 32*5 ), true),
						62 => (D_ipd(11)'last_event,  tpd_D_O((511 - 18)- 32*4 ), true),
						63 => (D_ipd(12)'last_event,  tpd_D_O((511 - 18)- 32*3 ), true),
						64=> (D_ipd(13)'last_event,  tpd_D_O((511 - 18)- 32*2 ), true),
						65=> (D_ipd(14)'last_event,  tpd_D_O((511 - 18)- 32*1 ), true), 
						66=> (D_ipd(15)'last_event,  tpd_D_O((511 - 18)- 32*0 ), true),
						67=> (CI_ipd'last_event, tpd_CI_O(13), true)  ,  
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(13), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(13),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(13),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(13),true)),
      Mode          => VitalTransport,
	  IgnoreDefaultDelay => TRUE,
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);  
	  
	  
	  	  	   VitalPathDelay01 (
      OutSignal     => O(14),
      GlitchData    => O_GlitchData(14),
      OutSignalName => "O(14)",
      OutTemp       => O_zd(14),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(14), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(14), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(14), true),
							3 => (A_ipd(0)'last_event,  tpd_A_O((511 - 17)- 32*15 ), true),
						4 => (A_ipd(1)'last_event,  tpd_A_O((511 - 17)- 32*14 ), true),
						5 => (A_ipd(2)'last_event,  tpd_A_O((511 - 17)- 32*13 ), true),
						6 => (A_ipd(3)'last_event,  tpd_A_O((511 - 17)- 32*12 ), true),
						7 => (A_ipd(4)'last_event,  tpd_A_O((511 - 17)- 32*11 ), true), 
						8 => (A_ipd(5)'last_event,  tpd_A_O((511 - 17)- 32*10 ), true),
						9 => (A_ipd(6)'last_event,  tpd_A_O((511 - 17)- 32*9 ), true),
						10 => (A_ipd(7)'last_event,  tpd_A_O((511 - 17)- 32*8 ), true),
						11=> (A_ipd(8)'last_event,  tpd_A_O((511 - 17)- 32*7 ), true),
						12 => (A_ipd(9)'last_event,  tpd_A_O((511 - 17)- 32*6 ), true),
						13 => (A_ipd(10)'last_event,  tpd_A_O((511 - 17)- 32*5 ), true),
						14 => (A_ipd(11)'last_event,  tpd_A_O((511 - 17)- 32*4 ), true),
						15 => (A_ipd(12)'last_event,  tpd_A_O((511 - 17)- 32*3 ), true),
						16=> (A_ipd(13)'last_event,  tpd_A_O((511 - 17)- 32*2), true),
						17=> (A_ipd(14)'last_event,  tpd_A_O((511 - 17)- 32*1 ), true), 
						18=> (A_ipd(15)'last_event,  tpd_A_O((511 - 17)- 32*0 ), true), 
						19=> (B_ipd(0)'last_event,  tpd_B_O((511 - 17)- 32*15 ), true),
						20 => (B_ipd(1)'last_event,  tpd_B_O((511 - 17)- 32*14 ), true),
						21 => (B_ipd(2)'last_event,  tpd_B_O((511 - 17)- 32*13 ), true),
						22 => (B_ipd(3)'last_event,  tpd_B_O((511 - 17)- 32*12 ), true),
						23=> (B_ipd(4)'last_event,  tpd_B_O((511 - 17)- 32*11 ), true), 
						24=> (B_ipd(5)'last_event,  tpd_B_O((511 - 17)- 32*10 ), true),
						25 => (B_ipd(6)'last_event,  tpd_B_O((511 - 17)- 32*9 ), true),
						26 => (B_ipd(7)'last_event,  tpd_B_O((511 - 17)- 32*8 ), true),
						27=> (B_ipd(8)'last_event,  tpd_B_O((511 - 17)- 32*7), true),
						28 => (B_ipd(9)'last_event,  tpd_B_O((511 - 17)- 32*6 ), true),
						29=> (B_ipd(10)'last_event,  tpd_B_O((511 - 17)- 32*5 ), true),
						30 => (B_ipd(11)'last_event,  tpd_B_O((511 - 17)- 32*4 ), true),
						31 => (B_ipd(12)'last_event,  tpd_B_O((511 - 17)- 32*3 ), true),
						32=> (B_ipd(13)'last_event,  tpd_B_O((511 - 17)- 32*2 ), true),
						33=> (B_ipd(14)'last_event,  tpd_B_O((511 - 17)- 32*1 ), true), 
						34=> (B_ipd(15)'last_event,  tpd_B_O((511 - 17)- 32*0 ), true),
						35=> (C_ipd(0)'last_event,  tpd_C_O((511 - 17)- 32*15 ), true),
						36 => (C_ipd(1)'last_event,  tpd_C_O((511 - 17)- 32*14 ), true),
						37 => (C_ipd(2)'last_event,  tpd_C_O((511 - 17)- 32*13 ), true),
						38 => (C_ipd(3)'last_event,  tpd_C_O((511 - 17)- 32*12 ), true),
						39=> (C_ipd(4)'last_event,  tpd_C_O((511 - 17)- 32*11 ), true), 
						40=> (C_ipd(5)'last_event,  tpd_C_O((511 - 17)- 32*10 ), true),
						41 => (C_ipd(6)'last_event,  tpd_C_O((511 - 17)- 32*9 ), true),
						42 => (C_ipd(7)'last_event,  tpd_C_O((511 - 17)- 32*8 ), true),
						43=> (C_ipd(8)'last_event,  tpd_C_O((511 - 17)- 32*7), true),
						44 => (C_ipd(9)'last_event,  tpd_C_O((511 - 17)- 32*6 ), true),
						45=> (C_ipd(10)'last_event,  tpd_C_O((511 - 17)- 32*5 ), true),
						46 => (C_ipd(11)'last_event,  tpd_C_O((511 - 17)- 32*4 ), true),
						47 => (C_ipd(12)'last_event,  tpd_C_O((511 - 17)- 32*3 ), true),
						48=> (C_ipd(13)'last_event,  tpd_C_O((511 - 17)- 32*2 ), true),
						49=> (C_ipd(14)'last_event,  tpd_C_O((511 - 17)- 32*1 ), true), 
						50=> (C_ipd(15)'last_event,  tpd_C_O((511 - 17)- 32*0 ), true),
						51=> (D_ipd(0)'last_event,  tpd_D_O((511 - 17)- 32*15 ), true),
						52 => (D_ipd(1)'last_event,  tpd_D_O((511 - 17)- 32*14 ), true),
						53 => (D_ipd(2)'last_event,  tpd_D_O((511 - 17)- 32*13 ), true),
						54 => (D_ipd(3)'last_event,  tpd_D_O((511 - 17)- 32*12 ), true),
						55=> (D_ipd(4)'last_event,  tpd_D_O((511 - 17)- 32*11 ), true), 
						56=> (D_ipd(5)'last_event,  tpd_D_O((511 - 17)- 32*10 ), true),
						57 => (D_ipd(6)'last_event,  tpd_D_O((511 - 17)- 32*9 ), true),
						58 => (D_ipd(7)'last_event,  tpd_D_O((511 - 17)- 32*8 ), true),
						59=> (D_ipd(8)'last_event,  tpd_D_O((511 - 17)- 32*7 ), true),
						60 => (D_ipd(9)'last_event,  tpd_D_O((511 - 17)- 32*6 ), true),
						61=> (D_ipd(10)'last_event,  tpd_D_O((511 - 17)- 32*5 ), true),
						62 => (D_ipd(11)'last_event,  tpd_D_O((511 - 17)- 32*4 ), true),
						63 => (D_ipd(12)'last_event,  tpd_D_O((511 - 17)- 32*3 ), true),
						64=> (D_ipd(13)'last_event,  tpd_D_O((511 - 17)- 32*2 ), true),
						65=> (D_ipd(14)'last_event,  tpd_D_O((511 - 17)- 32*1 ), true), 
						66=> (D_ipd(15)'last_event,  tpd_D_O((511 - 17)- 32*0 ), true),
						67=> (CI_ipd'last_event, tpd_CI_O(14), true)  ,  
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(14), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(14),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(14),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(14),true)),
      Mode          => VitalTransport,	   
	  IgnoreDefaultDelay => TRUE,
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);   
	  
	  
	  
	  	  	   VitalPathDelay01 (
      OutSignal     => O(15),
      GlitchData    => O_GlitchData(15),
      OutSignalName => "O(15)",
      OutTemp       => O_zd(15),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(15), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(15), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(15), true),
							3 => (A_ipd(0)'last_event,  tpd_A_O((511 - 16)- 32*15 ), true),
						4 => (A_ipd(1)'last_event,  tpd_A_O((511 - 16)- 32*14 ), true),
						5 => (A_ipd(2)'last_event,  tpd_A_O((511 - 16)- 32*13 ), true),
						6 => (A_ipd(3)'last_event,  tpd_A_O((511 - 16)- 32*12 ), true),
						7 => (A_ipd(4)'last_event,  tpd_A_O((511 - 16)- 32*11 ), true), 
						8 => (A_ipd(5)'last_event,  tpd_A_O((511 - 16)- 32*10 ), true),
						9 => (A_ipd(6)'last_event,  tpd_A_O((511 - 16)- 32*9 ), true),
						10 => (A_ipd(7)'last_event,  tpd_A_O((511 - 16)- 32*8 ), true),
						11=> (A_ipd(8)'last_event,  tpd_A_O((511 - 16)- 32*7 ), true),
						12 => (A_ipd(9)'last_event,  tpd_A_O((511 - 16)- 32*6 ), true),
						13 => (A_ipd(10)'last_event,  tpd_A_O((511 - 16)- 32*5 ), true),
						14 => (A_ipd(11)'last_event,  tpd_A_O((511 - 16)- 32*4 ), true),
						15 => (A_ipd(12)'last_event,  tpd_A_O((511 - 16)- 32*3 ), true),
						16=> (A_ipd(13)'last_event,  tpd_A_O((511 - 16)- 32*2), true),
						17=> (A_ipd(14)'last_event,  tpd_A_O((511 - 16)- 32*1 ), true), 
						18=> (A_ipd(15)'last_event,  tpd_A_O((511 - 16)- 32*0 ), true), 
						19=> (B_ipd(0)'last_event,  tpd_B_O((511 - 16)- 32*15 ), true),
						20 => (B_ipd(1)'last_event,  tpd_B_O((511 - 16)- 32*14 ), true),
						21 => (B_ipd(2)'last_event,  tpd_B_O((511 - 16)- 32*13 ), true),
						22 => (B_ipd(3)'last_event,  tpd_B_O((511 - 16)- 32*12 ), true),
						23=> (B_ipd(4)'last_event,  tpd_B_O((511 - 16)- 32*11 ), true), 
						24=> (B_ipd(5)'last_event,  tpd_B_O((511 - 16)- 32*10 ), true),
						25 => (B_ipd(6)'last_event,  tpd_B_O((511 - 16)- 32*9 ), true),
						26 => (B_ipd(7)'last_event,  tpd_B_O((511 - 16)- 32*8 ), true),
						27=> (B_ipd(8)'last_event,  tpd_B_O((511 - 16)- 32*7), true),
						28 => (B_ipd(9)'last_event,  tpd_B_O((511 - 16)- 32*6 ), true),
						29=> (B_ipd(10)'last_event,  tpd_B_O((511 - 16)- 32*5 ), true),
						30 => (B_ipd(11)'last_event,  tpd_B_O((511 - 16)- 32*4 ), true),
						31 => (B_ipd(12)'last_event,  tpd_B_O((511 - 16)- 32*3 ), true),
						32=> (B_ipd(13)'last_event,  tpd_B_O((511 - 16)- 32*2 ), true),
						33=> (B_ipd(14)'last_event,  tpd_B_O((511 - 16)- 32*1 ), true), 
						34=> (B_ipd(15)'last_event,  tpd_B_O((511 - 16)- 32*0 ), true),
						35=> (C_ipd(0)'last_event,  tpd_C_O((511 - 16)- 32*15 ), true),
						36 => (C_ipd(1)'last_event,  tpd_C_O((511 - 16)- 32*14 ), true),
						37 => (C_ipd(2)'last_event,  tpd_C_O((511 - 16)- 32*13 ), true),
						38 => (C_ipd(3)'last_event,  tpd_C_O((511 - 16)- 32*12 ), true),
						39=> (C_ipd(4)'last_event,  tpd_C_O((511 - 16)- 32*11 ), true), 
						40=> (C_ipd(5)'last_event,  tpd_C_O((511 - 16)- 32*10 ), true),
						41 => (C_ipd(6)'last_event,  tpd_C_O((511 - 16)- 32*9 ), true),
						42 => (C_ipd(7)'last_event,  tpd_C_O((511 - 16)- 32*8 ), true),
						43=> (C_ipd(8)'last_event,  tpd_C_O((511 - 16)- 32*7), true),
						44 => (C_ipd(9)'last_event,  tpd_C_O((511 - 16)- 32*6 ), true),
						45=> (C_ipd(10)'last_event,  tpd_C_O((511 - 16)- 32*5 ), true),
						46 => (C_ipd(11)'last_event,  tpd_C_O((511 - 16)- 32*4 ), true),
						47 => (C_ipd(12)'last_event,  tpd_C_O((511 - 16)- 32*3 ), true),
						48=> (C_ipd(13)'last_event,  tpd_C_O((511 - 16)- 32*2 ), true),
						49=> (C_ipd(14)'last_event,  tpd_C_O((511 - 16)- 32*1 ), true), 
						50=> (C_ipd(15)'last_event,  tpd_C_O((511 - 16)- 32*0 ), true),
						51=> (D_ipd(0)'last_event,  tpd_D_O((511 - 16)- 32*15 ), true),
						52 => (D_ipd(1)'last_event,  tpd_D_O((511 - 16)- 32*14 ), true),
						53 => (D_ipd(2)'last_event,  tpd_D_O((511 - 16)- 32*13 ), true),
						54 => (D_ipd(3)'last_event,  tpd_D_O((511 - 16)- 32*12 ), true),
						55=> (D_ipd(4)'last_event,  tpd_D_O((511 - 16)- 32*11 ), true), 
						56=> (D_ipd(5)'last_event,  tpd_D_O((511 - 16)- 32*10 ), true),
						57 => (D_ipd(6)'last_event,  tpd_D_O((511 - 16)- 32*9 ), true),
						58 => (D_ipd(7)'last_event,  tpd_D_O((511 - 16)- 32*8 ), true),
						59=> (D_ipd(8)'last_event,  tpd_D_O((511 - 16)- 32*7 ), true),
						60 => (D_ipd(9)'last_event,  tpd_D_O((511 - 16)- 32*6 ), true),
						61=> (D_ipd(10)'last_event,  tpd_D_O((511 - 16)- 32*5 ), true),
						62 => (D_ipd(11)'last_event,  tpd_D_O((511 - 16)- 32*4 ), true),
						63 => (D_ipd(12)'last_event,  tpd_D_O((511 - 16)- 32*3 ), true),
						64=> (D_ipd(13)'last_event,  tpd_D_O((511 - 16)- 32*2 ), true),
						65=> (D_ipd(14)'last_event,  tpd_D_O((511 - 16)- 32*1 ), true), 
						66=> (D_ipd(15)'last_event,  tpd_D_O((511 - 16)- 32*0 ), true),
						67=> (CI_ipd'last_event, tpd_CI_O(15), true)  ,  
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(15), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(15),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(15),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(15),true)),
      Mode          => VitalTransport,	 
	  IgnoreDefaultDelay => TRUE,  
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);	   
	  
	  
	  	  	   VitalPathDelay01 (
      OutSignal     => O(16),
      GlitchData    => O_GlitchData(16),
      OutSignalName => "O(16)",
      OutTemp       => O_zd(16),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(16), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(16), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(16), true),
							3 => (A_ipd(0)'last_event,  tpd_A_O((511 - 15)- 32*15 ), true),
						4 => (A_ipd(1)'last_event,  tpd_A_O((511 - 15)- 32*14 ), true),
						5 => (A_ipd(2)'last_event,  tpd_A_O((511 - 15)- 32*13 ), true),
						6 => (A_ipd(3)'last_event,  tpd_A_O((511 - 15)- 32*12 ), true),
						7 => (A_ipd(4)'last_event,  tpd_A_O((511 - 15)- 32*11 ), true), 
						8 => (A_ipd(5)'last_event,  tpd_A_O((511 - 15)- 32*10 ), true),
						9 => (A_ipd(6)'last_event,  tpd_A_O((511 - 15)- 32*9 ), true),
						10 => (A_ipd(7)'last_event,  tpd_A_O((511 - 15)- 32*8 ), true),
						11=> (A_ipd(8)'last_event,  tpd_A_O((511 - 15)- 32*7 ), true),
						12 => (A_ipd(9)'last_event,  tpd_A_O((511 - 15)- 32*6 ), true),
						13 => (A_ipd(10)'last_event,  tpd_A_O((511 - 15)- 32*5 ), true),
						14 => (A_ipd(11)'last_event,  tpd_A_O((511 - 15)- 32*4 ), true),
						15 => (A_ipd(12)'last_event,  tpd_A_O((511 - 15)- 32*3 ), true),
						16=> (A_ipd(13)'last_event,  tpd_A_O((511 - 15)- 32*2), true),
						17=> (A_ipd(14)'last_event,  tpd_A_O((511 - 15)- 32*1 ), true), 
						18=> (A_ipd(15)'last_event,  tpd_A_O((511 - 15)- 32*0 ), true), 
						19=> (B_ipd(0)'last_event,  tpd_B_O((511 - 15)- 32*15 ), true),
						20 => (B_ipd(1)'last_event,  tpd_B_O((511 - 15)- 32*14 ), true),
						21 => (B_ipd(2)'last_event,  tpd_B_O((511 - 15)- 32*13 ), true),
						22 => (B_ipd(3)'last_event,  tpd_B_O((511 - 15)- 32*12 ), true),
						23=> (B_ipd(4)'last_event,  tpd_B_O((511 - 15)- 32*11 ), true), 
						24=> (B_ipd(5)'last_event,  tpd_B_O((511 - 15)- 32*10 ), true),
						25 => (B_ipd(6)'last_event,  tpd_B_O((511 - 15)- 32*9 ), true),
						26 => (B_ipd(7)'last_event,  tpd_B_O((511 - 15)- 32*8 ), true),
						27=> (B_ipd(8)'last_event,  tpd_B_O((511 - 15)- 32*7), true),
						28 => (B_ipd(9)'last_event,  tpd_B_O((511 - 15)- 32*6 ), true),
						29=> (B_ipd(10)'last_event,  tpd_B_O((511 - 15)- 32*5 ), true),
						30 => (B_ipd(11)'last_event,  tpd_B_O((511 - 15)- 32*4 ), true),
						31 => (B_ipd(12)'last_event,  tpd_B_O((511 - 15)- 32*3 ), true),
						32=> (B_ipd(13)'last_event,  tpd_B_O((511 - 15)- 32*2 ), true),
						33=> (B_ipd(14)'last_event,  tpd_B_O((511 - 15)- 32*1 ), true), 
						34=> (B_ipd(15)'last_event,  tpd_B_O((511 - 15)- 32*0 ), true),
						35=> (C_ipd(0)'last_event,  tpd_C_O((511 - 15)- 32*15 ), true),
						36 => (C_ipd(1)'last_event,  tpd_C_O((511 - 15)- 32*14 ), true),
						37 => (C_ipd(2)'last_event,  tpd_C_O((511 - 15)- 32*13 ), true),
						38 => (C_ipd(3)'last_event,  tpd_C_O((511 - 15)- 32*12 ), true),
						39=> (C_ipd(4)'last_event,  tpd_C_O((511 - 15)- 32*11 ), true), 
						40=> (C_ipd(5)'last_event,  tpd_C_O((511 - 15)- 32*10 ), true),
						41 => (C_ipd(6)'last_event,  tpd_C_O((511 - 15)- 32*9 ), true),
						42 => (C_ipd(7)'last_event,  tpd_C_O((511 - 15)- 32*8 ), true),
						43=> (C_ipd(8)'last_event,  tpd_C_O((511 - 15)- 32*7), true),
						44 => (C_ipd(9)'last_event,  tpd_C_O((511 - 15)- 32*6 ), true),
						45=> (C_ipd(10)'last_event,  tpd_C_O((511 - 15)- 32*5 ), true),
						46 => (C_ipd(11)'last_event,  tpd_C_O((511 - 15)- 32*4 ), true),
						47 => (C_ipd(12)'last_event,  tpd_C_O((511 - 15)- 32*3 ), true),
						48=> (C_ipd(13)'last_event,  tpd_C_O((511 - 15)- 32*2 ), true),
						49=> (C_ipd(14)'last_event,  tpd_C_O((511 - 15)- 32*1 ), true), 
						50=> (C_ipd(15)'last_event,  tpd_C_O((511 - 15)- 32*0 ), true),
						51=> (D_ipd(0)'last_event,  tpd_D_O((511 - 15)- 32*15 ), true),
						52 => (D_ipd(1)'last_event,  tpd_D_O((511 - 15)- 32*14 ), true),
						53 => (D_ipd(2)'last_event,  tpd_D_O((511 - 15)- 32*13 ), true),
						54 => (D_ipd(3)'last_event,  tpd_D_O((511 - 15)- 32*12 ), true),
						55=> (D_ipd(4)'last_event,  tpd_D_O((511 - 15)- 32*11 ), true), 
						56=> (D_ipd(5)'last_event,  tpd_D_O((511 - 15)- 32*10 ), true),
						57 => (D_ipd(6)'last_event,  tpd_D_O((511 - 15)- 32*9 ), true),
						58 => (D_ipd(7)'last_event,  tpd_D_O((511 - 15)- 32*8 ), true),
						59=> (D_ipd(8)'last_event,  tpd_D_O((511 - 15)- 32*7 ), true),
						60 => (D_ipd(9)'last_event,  tpd_D_O((511 - 15)- 32*6 ), true),
						61=> (D_ipd(10)'last_event,  tpd_D_O((511 - 15)- 32*5 ), true),
						62 => (D_ipd(11)'last_event,  tpd_D_O((511 - 15)- 32*4 ), true),
						63 => (D_ipd(12)'last_event,  tpd_D_O((511 - 15)- 32*3 ), true),
						64=> (D_ipd(13)'last_event,  tpd_D_O((511 - 15)- 32*2 ), true),
						65=> (D_ipd(14)'last_event,  tpd_D_O((511 - 15)- 32*1 ), true), 
						66=> (D_ipd(15)'last_event,  tpd_D_O((511 - 15)- 32*0 ), true),
						67=> (CI_ipd'last_event, tpd_CI_O(16), true)  ,  
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(16), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(16),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(16),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(16),true)),
      Mode          => VitalTransport,	 
	  IgnoreDefaultDelay => TRUE,	
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);
	  
	  
	  	  	  	   VitalPathDelay01 (
      OutSignal     => O(17),
      GlitchData    => O_GlitchData(17),
      OutSignalName => "O(17)",
      OutTemp       => O_zd(17),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(17), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(17), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(17), true),
						3 => (A_ipd(0)'last_event,  tpd_A_O((511 - 14)- 32*15 ), true),
						4 => (A_ipd(1)'last_event,  tpd_A_O((511 - 14)- 32*14 ), true),
						5 => (A_ipd(2)'last_event,  tpd_A_O((511 - 14)- 32*13 ), true),
						6 => (A_ipd(3)'last_event,  tpd_A_O((511 - 14)- 32*12 ), true),
						7 => (A_ipd(4)'last_event,  tpd_A_O((511 - 14)- 32*11 ), true), 
						8 => (A_ipd(5)'last_event,  tpd_A_O((511 - 14)- 32*10 ), true),
						9 => (A_ipd(6)'last_event,  tpd_A_O((511 - 14)- 32*9 ), true),
						10 => (A_ipd(7)'last_event,  tpd_A_O((511 - 14)- 32*8 ), true),
						11=> (A_ipd(8)'last_event,  tpd_A_O((511 - 14)- 32*7 ), true),
						12 => (A_ipd(9)'last_event,  tpd_A_O((511 - 14)- 32*6 ), true),
						13 => (A_ipd(10)'last_event,  tpd_A_O((511 - 14)- 32*5 ), true),
						14 => (A_ipd(11)'last_event,  tpd_A_O((511 - 14)- 32*4 ), true),
						15 => (A_ipd(12)'last_event,  tpd_A_O((511 - 14)- 32*3 ), true),
						16=> (A_ipd(13)'last_event,  tpd_A_O((511 - 14)- 32*2), true),
						17=> (A_ipd(14)'last_event,  tpd_A_O((511 - 14)- 32*1 ), true), 
						18=> (A_ipd(15)'last_event,  tpd_A_O((511 - 14)- 32*0 ), true), 
						19=> (B_ipd(0)'last_event,  tpd_B_O((511 - 14)- 32*15 ), true),
						20 => (B_ipd(1)'last_event,  tpd_B_O((511 - 14)- 32*14 ), true),
						21 => (B_ipd(2)'last_event,  tpd_B_O((511 - 14)- 32*13 ), true),
						22 => (B_ipd(3)'last_event,  tpd_B_O((511 - 14)- 32*12 ), true),
						23=> (B_ipd(4)'last_event,  tpd_B_O((511 - 14)- 32*11 ), true), 
						24=> (B_ipd(5)'last_event,  tpd_B_O((511 - 14)- 32*10 ), true),
						25 => (B_ipd(6)'last_event,  tpd_B_O((511 - 14)- 32*9 ), true),
						26 => (B_ipd(7)'last_event,  tpd_B_O((511 - 14)- 32*8 ), true),
						27=> (B_ipd(8)'last_event,  tpd_B_O((511 - 14)- 32*7), true),
						28 => (B_ipd(9)'last_event,  tpd_B_O((511 - 14)- 32*6 ), true),
						29=> (B_ipd(10)'last_event,  tpd_B_O((511 - 14)- 32*5 ), true),
						30 => (B_ipd(11)'last_event,  tpd_B_O((511 - 14)- 32*4 ), true),
						31 => (B_ipd(12)'last_event,  tpd_B_O((511 - 14)- 32*3 ), true),
						32=> (B_ipd(13)'last_event,  tpd_B_O((511 - 14)- 32*2 ), true),
						33=> (B_ipd(14)'last_event,  tpd_B_O((511 - 14)- 32*1 ), true), 
						34=> (B_ipd(15)'last_event,  tpd_B_O((511 - 14)- 32*0 ), true),
						35=> (C_ipd(0)'last_event,  tpd_C_O((511 - 14)- 32*15 ), true),
						36 => (C_ipd(1)'last_event,  tpd_C_O((511 - 14)- 32*14 ), true),
						37 => (C_ipd(2)'last_event,  tpd_C_O((511 - 14)- 32*13 ), true),
						38 => (C_ipd(3)'last_event,  tpd_C_O((511 - 14)- 32*12 ), true),
						39=> (C_ipd(4)'last_event,  tpd_C_O((511 - 14)- 32*11 ), true), 
						40=> (C_ipd(5)'last_event,  tpd_C_O((511 - 14)- 32*10 ), true),
						41 => (C_ipd(6)'last_event,  tpd_C_O((511 - 14)- 32*9 ), true),
						42 => (C_ipd(7)'last_event,  tpd_C_O((511 - 14)- 32*8 ), true),
						43=> (C_ipd(8)'last_event,  tpd_C_O((511 - 14)- 32*7), true),
						44 => (C_ipd(9)'last_event,  tpd_C_O((511 - 14)- 32*6 ), true),
						45=> (C_ipd(10)'last_event,  tpd_C_O((511 - 14)- 32*5 ), true),
						46 => (C_ipd(11)'last_event,  tpd_C_O((511 - 14)- 32*4 ), true),
						47 => (C_ipd(12)'last_event,  tpd_C_O((511 - 14)- 32*3 ), true),
						48=> (C_ipd(13)'last_event,  tpd_C_O((511 - 14)- 32*2 ), true),
						49=> (C_ipd(14)'last_event,  tpd_C_O((511 - 14)- 32*1 ), true), 
						50=> (C_ipd(15)'last_event,  tpd_C_O((511 - 14)- 32*0 ), true),
						51=> (D_ipd(0)'last_event,  tpd_D_O((511 - 14)- 32*15 ), true),
						52 => (D_ipd(1)'last_event,  tpd_D_O((511 - 14)- 32*14 ), true),
						53 => (D_ipd(2)'last_event,  tpd_D_O((511 - 14)- 32*13 ), true),
						54 => (D_ipd(3)'last_event,  tpd_D_O((511 - 14)- 32*12 ), true),
						55=> (D_ipd(4)'last_event,  tpd_D_O((511 - 14)- 32*11 ), true), 
						56=> (D_ipd(5)'last_event,  tpd_D_O((511 - 14)- 32*10 ), true),
						57 => (D_ipd(6)'last_event,  tpd_D_O((511 - 14)- 32*9 ), true),
						58 => (D_ipd(7)'last_event,  tpd_D_O((511 - 14)- 32*8 ), true),
						59=> (D_ipd(8)'last_event,  tpd_D_O((511 - 14)- 32*7 ), true),
						60 => (D_ipd(9)'last_event,  tpd_D_O((511 - 14)- 32*6 ), true),
						61=> (D_ipd(10)'last_event,  tpd_D_O((511 - 14)- 32*5 ), true),
						62 => (D_ipd(11)'last_event,  tpd_D_O((511 - 14)- 32*4 ), true),
						63 => (D_ipd(12)'last_event,  tpd_D_O((511 - 14)- 32*3 ), true),
						64=> (D_ipd(13)'last_event,  tpd_D_O((511 - 14)- 32*2 ), true),
						65=> (D_ipd(14)'last_event,  tpd_D_O((511 - 14)- 32*1 ), true), 
						66=> (D_ipd(15)'last_event,  tpd_D_O((511 - 14)- 32*0 ), true),
						67=> (CI_ipd'last_event, tpd_CI_O(17), true)  ,  
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(17), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(17),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(17),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(17),true)),
      Mode          => VitalTransport,	   
	  IgnoreDefaultDelay => TRUE,
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);  
	  
	  
	  	  	  	   VitalPathDelay01 (
      OutSignal     => O(18),
      GlitchData    => O_GlitchData(18),
      OutSignalName => "O(18)",
      OutTemp       => O_zd(18),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(18), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(18), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(18), true),
							3 => (A_ipd(0)'last_event,  tpd_A_O((511 - 13)- 32*15 ), true),
						4 => (A_ipd(1)'last_event,  tpd_A_O((511 - 13)- 32*14 ), true),
						5 => (A_ipd(2)'last_event,  tpd_A_O((511 - 13)- 32*13 ), true),
						6 => (A_ipd(3)'last_event,  tpd_A_O((511 - 13)- 32*12 ), true),
						7 => (A_ipd(4)'last_event,  tpd_A_O((511 - 13)- 32*11 ), true), 
						8 => (A_ipd(5)'last_event,  tpd_A_O((511 - 13)- 32*10 ), true),
						9 => (A_ipd(6)'last_event,  tpd_A_O((511 - 13)- 32*9 ), true),
						10 => (A_ipd(7)'last_event,  tpd_A_O((511 - 13)- 32*8 ), true),
						11=> (A_ipd(8)'last_event,  tpd_A_O((511 - 13)- 32*7 ), true),
						12 => (A_ipd(9)'last_event,  tpd_A_O((511 - 13)- 32*6 ), true),
						13 => (A_ipd(10)'last_event,  tpd_A_O((511 - 13)- 32*5 ), true),
						14 => (A_ipd(11)'last_event,  tpd_A_O((511 - 13)- 32*4 ), true),
						15 => (A_ipd(12)'last_event,  tpd_A_O((511 - 13)- 32*3 ), true),
						16=> (A_ipd(13)'last_event,  tpd_A_O((511 - 13)- 32*2), true),
						17=> (A_ipd(14)'last_event,  tpd_A_O((511 - 13)- 32*1 ), true), 
						18=> (A_ipd(15)'last_event,  tpd_A_O((511 - 13)- 32*0 ), true), 
						19=> (B_ipd(0)'last_event,  tpd_B_O((511 - 13)- 32*15 ), true),
						20 => (B_ipd(1)'last_event,  tpd_B_O((511 - 13)- 32*14 ), true),
						21 => (B_ipd(2)'last_event,  tpd_B_O((511 - 13)- 32*13 ), true),
						22 => (B_ipd(3)'last_event,  tpd_B_O((511 - 13)- 32*12 ), true),
						23=> (B_ipd(4)'last_event,  tpd_B_O((511 - 13)- 32*11 ), true), 
						24=> (B_ipd(5)'last_event,  tpd_B_O((511 - 13)- 32*10 ), true),
						25 => (B_ipd(6)'last_event,  tpd_B_O((511 - 13)- 32*9 ), true),
						26 => (B_ipd(7)'last_event,  tpd_B_O((511 - 13)- 32*8 ), true),
						27=> (B_ipd(8)'last_event,  tpd_B_O((511 - 13)- 32*7), true),
						28 => (B_ipd(9)'last_event,  tpd_B_O((511 - 13)- 32*6 ), true),
						29=> (B_ipd(10)'last_event,  tpd_B_O((511 - 13)- 32*5 ), true),
						30 => (B_ipd(11)'last_event,  tpd_B_O((511 - 13)- 32*4 ), true),
						31 => (B_ipd(12)'last_event,  tpd_B_O((511 - 13)- 32*3 ), true),
						32=> (B_ipd(13)'last_event,  tpd_B_O((511 - 13)- 32*2 ), true),
						33=> (B_ipd(14)'last_event,  tpd_B_O((511 - 13)- 32*1 ), true), 
						34=> (B_ipd(15)'last_event,  tpd_B_O((511 - 13)- 32*0 ), true),
						35=> (C_ipd(0)'last_event,  tpd_C_O((511 - 13)- 32*15 ), true),
						36 => (C_ipd(1)'last_event,  tpd_C_O((511 - 13)- 32*14 ), true),
						37 => (C_ipd(2)'last_event,  tpd_C_O((511 - 13)- 32*13 ), true),
						38 => (C_ipd(3)'last_event,  tpd_C_O((511 - 13)- 32*12 ), true),
						39=> (C_ipd(4)'last_event,  tpd_C_O((511 - 13)- 32*11 ), true), 
						40=> (C_ipd(5)'last_event,  tpd_C_O((511 - 13)- 32*10 ), true),
						41 => (C_ipd(6)'last_event,  tpd_C_O((511 - 13)- 32*9 ), true),
						42 => (C_ipd(7)'last_event,  tpd_C_O((511 - 13)- 32*8 ), true),
						43=> (C_ipd(8)'last_event,  tpd_C_O((511 - 13)- 32*7), true),
						44 => (C_ipd(9)'last_event,  tpd_C_O((511 - 13)- 32*6 ), true),
						45=> (C_ipd(10)'last_event,  tpd_C_O((511 - 13)- 32*5 ), true),
						46 => (C_ipd(11)'last_event,  tpd_C_O((511 - 13)- 32*4 ), true),
						47 => (C_ipd(12)'last_event,  tpd_C_O((511 - 13)- 32*3 ), true),
						48=> (C_ipd(13)'last_event,  tpd_C_O((511 - 13)- 32*2 ), true),
						49=> (C_ipd(14)'last_event,  tpd_C_O((511 - 13)- 32*1 ), true), 
						50=> (C_ipd(15)'last_event,  tpd_C_O((511 - 13)- 32*0 ), true),
						51=> (D_ipd(0)'last_event,  tpd_D_O((511 - 13)- 32*15 ), true),
						52 => (D_ipd(1)'last_event,  tpd_D_O((511 - 13)- 32*14 ), true),
						53 => (D_ipd(2)'last_event,  tpd_D_O((511 - 13)- 32*13 ), true),
						54 => (D_ipd(3)'last_event,  tpd_D_O((511 - 13)- 32*12 ), true),
						55=> (D_ipd(4)'last_event,  tpd_D_O((511 - 13)- 32*11 ), true), 
						56=> (D_ipd(5)'last_event,  tpd_D_O((511 - 13)- 32*10 ), true),
						57 => (D_ipd(6)'last_event,  tpd_D_O((511 - 13)- 32*9 ), true),
						58 => (D_ipd(7)'last_event,  tpd_D_O((511 - 13)- 32*8 ), true),
						59=> (D_ipd(8)'last_event,  tpd_D_O((511 - 13)- 32*7 ), true),
						60 => (D_ipd(9)'last_event,  tpd_D_O((511 - 13)- 32*6 ), true),
						61=> (D_ipd(10)'last_event,  tpd_D_O((511 - 13)- 32*5 ), true),
						62 => (D_ipd(11)'last_event,  tpd_D_O((511 - 13)- 32*4 ), true),
						63 => (D_ipd(12)'last_event,  tpd_D_O((511 - 13)- 32*3 ), true),
						64=> (D_ipd(13)'last_event,  tpd_D_O((511 - 13)- 32*2 ), true),
						65=> (D_ipd(14)'last_event,  tpd_D_O((511 - 13)- 32*1 ), true), 
						66=> (D_ipd(15)'last_event,  tpd_D_O((511 - 13)- 32*0 ), true),
						67=> (CI_ipd'last_event, tpd_CI_O(18), true)  ,  
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(18), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(18),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(18),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(18),true)),
      Mode          => VitalTransport,
	  IgnoreDefaultDelay => TRUE, 
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);  
	  
	  
	  	  	  	   VitalPathDelay01 (
      OutSignal     => O(19),
      GlitchData    => O_GlitchData(19),
      OutSignalName => "O(19)",
      OutTemp       => O_zd(19),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(19), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(19), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(19), true),
							3 => (A_ipd(0)'last_event,  tpd_A_O((511 - 12)- 32*15 ), true),
						4 => (A_ipd(1)'last_event,  tpd_A_O((511 - 12)- 32*14 ), true),
						5 => (A_ipd(2)'last_event,  tpd_A_O((511 - 12)- 32*13 ), true),
						6 => (A_ipd(3)'last_event,  tpd_A_O((511 - 12)- 32*12 ), true),
						7 => (A_ipd(4)'last_event,  tpd_A_O((511 - 12)- 32*11 ), true), 
						8 => (A_ipd(5)'last_event,  tpd_A_O((511 - 12)- 32*10 ), true),
						9 => (A_ipd(6)'last_event,  tpd_A_O((511 - 12)- 32*9 ), true),
						10 => (A_ipd(7)'last_event,  tpd_A_O((511 - 12)- 32*8 ), true),
						11=> (A_ipd(8)'last_event,  tpd_A_O((511 - 12)- 32*7 ), true),
						12 => (A_ipd(9)'last_event,  tpd_A_O((511 - 12)- 32*6 ), true),
						13 => (A_ipd(10)'last_event,  tpd_A_O((511 - 12)- 32*5 ), true),
						14 => (A_ipd(11)'last_event,  tpd_A_O((511 - 12)- 32*4 ), true),
						15 => (A_ipd(12)'last_event,  tpd_A_O((511 - 12)- 32*3 ), true),
						16=> (A_ipd(13)'last_event,  tpd_A_O((511 - 12)- 32*2), true),
						17=> (A_ipd(14)'last_event,  tpd_A_O((511 - 12)- 32*1 ), true), 
						18=> (A_ipd(15)'last_event,  tpd_A_O((511 - 12)- 32*0 ), true), 
						19=> (B_ipd(0)'last_event,  tpd_B_O((511 - 12)- 32*15 ), true),
						20 => (B_ipd(1)'last_event,  tpd_B_O((511 - 12)- 32*14 ), true),
						21 => (B_ipd(2)'last_event,  tpd_B_O((511 - 12)- 32*13 ), true),
						22 => (B_ipd(3)'last_event,  tpd_B_O((511 - 12)- 32*12 ), true),
						23=> (B_ipd(4)'last_event,  tpd_B_O((511 - 12)- 32*11 ), true), 
						24=> (B_ipd(5)'last_event,  tpd_B_O((511 - 12)- 32*10 ), true),
						25 => (B_ipd(6)'last_event,  tpd_B_O((511 - 12)- 32*9 ), true),
						26 => (B_ipd(7)'last_event,  tpd_B_O((511 - 12)- 32*8 ), true),
						27=> (B_ipd(8)'last_event,  tpd_B_O((511 - 12)- 32*7), true),
						28 => (B_ipd(9)'last_event,  tpd_B_O((511 - 12)- 32*6 ), true),
						29=> (B_ipd(10)'last_event,  tpd_B_O((511 - 12)- 32*5 ), true),
						30 => (B_ipd(11)'last_event,  tpd_B_O((511 - 12)- 32*4 ), true),
						31 => (B_ipd(12)'last_event,  tpd_B_O((511 - 12)- 32*3 ), true),
						32=> (B_ipd(13)'last_event,  tpd_B_O((511 - 12)- 32*2 ), true),
						33=> (B_ipd(14)'last_event,  tpd_B_O((511 - 12)- 32*1 ), true), 
						34=> (B_ipd(15)'last_event,  tpd_B_O((511 - 12)- 32*0 ), true),
						35=> (C_ipd(0)'last_event,  tpd_C_O((511 - 12)- 32*15 ), true),
						36 => (C_ipd(1)'last_event,  tpd_C_O((511 - 12)- 32*14 ), true),
						37 => (C_ipd(2)'last_event,  tpd_C_O((511 - 12)- 32*13 ), true),
						38 => (C_ipd(3)'last_event,  tpd_C_O((511 - 12)- 32*12 ), true),
						39=> (C_ipd(4)'last_event,  tpd_C_O((511 - 12)- 32*11 ), true), 
						40=> (C_ipd(5)'last_event,  tpd_C_O((511 - 12)- 32*10 ), true),
						41 => (C_ipd(6)'last_event,  tpd_C_O((511 - 12)- 32*9 ), true),
						42 => (C_ipd(7)'last_event,  tpd_C_O((511 - 12)- 32*8 ), true),
						43=> (C_ipd(8)'last_event,  tpd_C_O((511 - 12)- 32*7), true),
						44 => (C_ipd(9)'last_event,  tpd_C_O((511 - 12)- 32*6 ), true),
						45=> (C_ipd(10)'last_event,  tpd_C_O((511 - 12)- 32*5 ), true),
						46 => (C_ipd(11)'last_event,  tpd_C_O((511 - 12)- 32*4 ), true),
						47 => (C_ipd(12)'last_event,  tpd_C_O((511 - 12)- 32*3 ), true),
						48=> (C_ipd(13)'last_event,  tpd_C_O((511 - 12)- 32*2 ), true),
						49=> (C_ipd(14)'last_event,  tpd_C_O((511 - 12)- 32*1 ), true), 
						50=> (C_ipd(15)'last_event,  tpd_C_O((511 - 12)- 32*0 ), true),
						51=> (D_ipd(0)'last_event,  tpd_D_O((511 - 12)- 32*15 ), true),
						52 => (D_ipd(1)'last_event,  tpd_D_O((511 - 12)- 32*14 ), true),
						53 => (D_ipd(2)'last_event,  tpd_D_O((511 - 12)- 32*13 ), true),
						54 => (D_ipd(3)'last_event,  tpd_D_O((511 - 12)- 32*12 ), true),
						55=> (D_ipd(4)'last_event,  tpd_D_O((511 - 12)- 32*11 ), true), 
						56=> (D_ipd(5)'last_event,  tpd_D_O((511 - 12)- 32*10 ), true),
						57 => (D_ipd(6)'last_event,  tpd_D_O((511 - 12)- 32*9 ), true),
						58 => (D_ipd(7)'last_event,  tpd_D_O((511 - 12)- 32*8 ), true),
						59=> (D_ipd(8)'last_event,  tpd_D_O((511 - 12)- 32*7 ), true),
						60 => (D_ipd(9)'last_event,  tpd_D_O((511 - 12)- 32*6 ), true),
						61=> (D_ipd(10)'last_event,  tpd_D_O((511 - 12)- 32*5 ), true),
						62 => (D_ipd(11)'last_event,  tpd_D_O((511 - 12)- 32*4 ), true),
						63 => (D_ipd(12)'last_event,  tpd_D_O((511 - 12)- 32*3 ), true),
						64=> (D_ipd(13)'last_event,  tpd_D_O((511 - 12)- 32*2 ), true),
						65=> (D_ipd(14)'last_event,  tpd_D_O((511 - 12)- 32*1 ), true), 
						66=> (D_ipd(15)'last_event,  tpd_D_O((511 - 12)- 32*0 ), true),
						67=> (CI_ipd'last_event, tpd_CI_O(19), true)  ,  
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(19), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(19),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(19),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(19),true)),
      Mode          => VitalTransport,	
	  IgnoreDefaultDelay => TRUE, 
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);  
	  
	  
	  
	  	  	  	   VitalPathDelay01 (
      OutSignal     => O(20),
      GlitchData    => O_GlitchData(20),
      OutSignalName => "O(20)",
      OutTemp       => O_zd(20),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(20), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(20), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(20), true),
						3 => (A_ipd(0)'last_event,  tpd_A_O((511 - 11)- 32*15 ), true),
						4 => (A_ipd(1)'last_event,  tpd_A_O((511 - 11)- 32*14 ), true),
						5 => (A_ipd(2)'last_event,  tpd_A_O((511 - 11)- 32*13 ), true),
						6 => (A_ipd(3)'last_event,  tpd_A_O((511 - 11)- 32*12 ), true),
						7 => (A_ipd(4)'last_event,  tpd_A_O((511 - 11)- 32*11 ), true), 
						8 => (A_ipd(5)'last_event,  tpd_A_O((511 - 11)- 32*10 ), true),
						9 => (A_ipd(6)'last_event,  tpd_A_O((511 - 11)- 32*9 ), true),
						10 => (A_ipd(7)'last_event,  tpd_A_O((511 - 11)- 32*8 ), true),
						11=> (A_ipd(8)'last_event,  tpd_A_O((511 - 11)- 32*7 ), true),
						12 => (A_ipd(9)'last_event,  tpd_A_O((511 - 11)- 32*6 ), true),
						13 => (A_ipd(10)'last_event,  tpd_A_O((511 - 11)- 32*5 ), true),
						14 => (A_ipd(11)'last_event,  tpd_A_O((511 - 11)- 32*4 ), true),
						15 => (A_ipd(12)'last_event,  tpd_A_O((511 - 11)- 32*3 ), true),
						16=> (A_ipd(13)'last_event,  tpd_A_O((511 - 11)- 32*2), true),
						17=> (A_ipd(14)'last_event,  tpd_A_O((511 - 11)- 32*1 ), true), 
						18=> (A_ipd(15)'last_event,  tpd_A_O((511 - 11)- 32*0 ), true), 
						19=> (B_ipd(0)'last_event,  tpd_B_O((511 - 11)- 32*15 ), true),
						20 => (B_ipd(1)'last_event,  tpd_B_O((511 - 11)- 32*14 ), true),
						21 => (B_ipd(2)'last_event,  tpd_B_O((511 - 11)- 32*13 ), true),
						22 => (B_ipd(3)'last_event,  tpd_B_O((511 - 11)- 32*12 ), true),
						23=> (B_ipd(4)'last_event,  tpd_B_O((511 - 11)- 32*11 ), true), 
						24=> (B_ipd(5)'last_event,  tpd_B_O((511 - 11)- 32*10 ), true),
						25 => (B_ipd(6)'last_event,  tpd_B_O((511 - 11)- 32*9 ), true),
						26 => (B_ipd(7)'last_event,  tpd_B_O((511 - 11)- 32*8 ), true),
						27=> (B_ipd(8)'last_event,  tpd_B_O((511 - 11)- 32*7), true),
						28 => (B_ipd(9)'last_event,  tpd_B_O((511 - 11)- 32*6 ), true),
						29=> (B_ipd(10)'last_event,  tpd_B_O((511 - 11)- 32*5 ), true),
						30 => (B_ipd(11)'last_event,  tpd_B_O((511 - 11)- 32*4 ), true),
						31 => (B_ipd(12)'last_event,  tpd_B_O((511 - 11)- 32*3 ), true),
						32=> (B_ipd(13)'last_event,  tpd_B_O((511 - 11)- 32*2 ), true),
						33=> (B_ipd(14)'last_event,  tpd_B_O((511 - 11)- 32*1 ), true), 
						34=> (B_ipd(15)'last_event,  tpd_B_O((511 - 11)- 32*0 ), true),
						35=> (C_ipd(0)'last_event,  tpd_C_O((511 - 11)- 32*15 ), true),
						36 => (C_ipd(1)'last_event,  tpd_C_O((511 - 11)- 32*14 ), true),
						37 => (C_ipd(2)'last_event,  tpd_C_O((511 - 11)- 32*13 ), true),
						38 => (C_ipd(3)'last_event,  tpd_C_O((511 - 11)- 32*12 ), true),
						39=> (C_ipd(4)'last_event,  tpd_C_O((511 - 11)- 32*11 ), true), 
						40=> (C_ipd(5)'last_event,  tpd_C_O((511 - 11)- 32*10 ), true),
						41 => (C_ipd(6)'last_event,  tpd_C_O((511 - 11)- 32*9 ), true),
						42 => (C_ipd(7)'last_event,  tpd_C_O((511 - 11)- 32*8 ), true),
						43=> (C_ipd(8)'last_event,  tpd_C_O((511 - 11)- 32*7), true),
						44 => (C_ipd(9)'last_event,  tpd_C_O((511 - 11)- 32*6 ), true),
						45=> (C_ipd(10)'last_event,  tpd_C_O((511 - 11)- 32*5 ), true),
						46 => (C_ipd(11)'last_event,  tpd_C_O((511 - 11)- 32*4 ), true),
						47 => (C_ipd(12)'last_event,  tpd_C_O((511 - 11)- 32*3 ), true),
						48=> (C_ipd(13)'last_event,  tpd_C_O((511 - 11)- 32*2 ), true),
						49=> (C_ipd(14)'last_event,  tpd_C_O((511 - 11)- 32*1 ), true), 
						50=> (C_ipd(15)'last_event,  tpd_C_O((511 - 11)- 32*0 ), true),
						51=> (D_ipd(0)'last_event,  tpd_D_O((511 - 11)- 32*15 ), true),
						52 => (D_ipd(1)'last_event,  tpd_D_O((511 - 11)- 32*14 ), true),
						53 => (D_ipd(2)'last_event,  tpd_D_O((511 - 11)- 32*13 ), true),
						54 => (D_ipd(3)'last_event,  tpd_D_O((511 - 11)- 32*12 ), true),
						55=> (D_ipd(4)'last_event,  tpd_D_O((511 - 11)- 32*11 ), true), 
						56=> (D_ipd(5)'last_event,  tpd_D_O((511 - 11)- 32*10 ), true),
						57 => (D_ipd(6)'last_event,  tpd_D_O((511 - 11)- 32*9 ), true),
						58 => (D_ipd(7)'last_event,  tpd_D_O((511 - 11)- 32*8 ), true),
						59=> (D_ipd(8)'last_event,  tpd_D_O((511 - 11)- 32*7 ), true),
						60 => (D_ipd(9)'last_event,  tpd_D_O((511 - 11)- 32*6 ), true),
						61=> (D_ipd(10)'last_event,  tpd_D_O((511 - 11)- 32*5 ), true),
						62 => (D_ipd(11)'last_event,  tpd_D_O((511 - 11)- 32*4 ), true),
						63 => (D_ipd(12)'last_event,  tpd_D_O((511 - 11)- 32*3 ), true),
						64=> (D_ipd(13)'last_event,  tpd_D_O((511 - 11)- 32*2 ), true),
						65=> (D_ipd(14)'last_event,  tpd_D_O((511 - 11)- 32*1 ), true), 
						66=> (D_ipd(15)'last_event,  tpd_D_O((511 - 11)- 32*0 ), true),
						67=> (CI_ipd'last_event, tpd_CI_O(20), true)  ,  
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(20), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(20),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(20),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(20),true)),
      Mode          => VitalTransport,	
	  IgnoreDefaultDelay => TRUE,
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);  
	  
	  
	  
	  	  	  	   VitalPathDelay01 (
      OutSignal     => O(21),
      GlitchData    => O_GlitchData(21),
      OutSignalName => "O(21)",
      OutTemp       => O_zd(21),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(21), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(21), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(21), true),
							3 => (A_ipd(0)'last_event,  tpd_A_O((511 - 10)- 32*15 ), true),
						4 => (A_ipd(1)'last_event,  tpd_A_O((511 - 10)- 32*14 ), true),
						5 => (A_ipd(2)'last_event,  tpd_A_O((511 - 10)- 32*13 ), true),
						6 => (A_ipd(3)'last_event,  tpd_A_O((511 - 10)- 32*12 ), true),
						7 => (A_ipd(4)'last_event,  tpd_A_O((511 - 10)- 32*11 ), true), 
						8 => (A_ipd(5)'last_event,  tpd_A_O((511 - 10)- 32*10 ), true),
						9 => (A_ipd(6)'last_event,  tpd_A_O((511 - 10)- 32*9 ), true),
						10 => (A_ipd(7)'last_event,  tpd_A_O((511 - 10)- 32*8 ), true),
						11=> (A_ipd(8)'last_event,  tpd_A_O((511 - 10)- 32*7 ), true),
						12 => (A_ipd(9)'last_event,  tpd_A_O((511 - 10)- 32*6 ), true),
						13 => (A_ipd(10)'last_event,  tpd_A_O((511 - 10)- 32*5 ), true),
						14 => (A_ipd(11)'last_event,  tpd_A_O((511 - 10)- 32*4 ), true),
						15 => (A_ipd(12)'last_event,  tpd_A_O((511 - 10)- 32*3 ), true),
						16=> (A_ipd(13)'last_event,  tpd_A_O((511 - 10)- 32*2), true),
						17=> (A_ipd(14)'last_event,  tpd_A_O((511 - 10)- 32*1 ), true), 
						18=> (A_ipd(15)'last_event,  tpd_A_O((511 - 10)- 32*0 ), true), 
						19=> (B_ipd(0)'last_event,  tpd_B_O((511 - 10)- 32*15 ), true),
						20 => (B_ipd(1)'last_event,  tpd_B_O((511 - 10)- 32*14 ), true),
						21 => (B_ipd(2)'last_event,  tpd_B_O((511 - 10)- 32*13 ), true),
						22 => (B_ipd(3)'last_event,  tpd_B_O((511 - 10)- 32*12 ), true),
						23=> (B_ipd(4)'last_event,  tpd_B_O((511 - 10)- 32*11 ), true), 
						24=> (B_ipd(5)'last_event,  tpd_B_O((511 - 10)- 32*10 ), true),
						25 => (B_ipd(6)'last_event,  tpd_B_O((511 - 10)- 32*9 ), true),
						26 => (B_ipd(7)'last_event,  tpd_B_O((511 - 10)- 32*8 ), true),
						27=> (B_ipd(8)'last_event,  tpd_B_O((511 - 10)- 32*7), true),
						28 => (B_ipd(9)'last_event,  tpd_B_O((511 - 10)- 32*6 ), true),
						29=> (B_ipd(10)'last_event,  tpd_B_O((511 - 10)- 32*5 ), true),
						30 => (B_ipd(11)'last_event,  tpd_B_O((511 - 10)- 32*4 ), true),
						31 => (B_ipd(12)'last_event,  tpd_B_O((511 - 10)- 32*3 ), true),
						32=> (B_ipd(13)'last_event,  tpd_B_O((511 - 10)- 32*2 ), true),
						33=> (B_ipd(14)'last_event,  tpd_B_O((511 - 10)- 32*1 ), true), 
						34=> (B_ipd(15)'last_event,  tpd_B_O((511 - 10)- 32*0 ), true),
						35=> (C_ipd(0)'last_event,  tpd_C_O((511 - 10)- 32*15 ), true),
						36 => (C_ipd(1)'last_event,  tpd_C_O((511 - 10)- 32*14 ), true),
						37 => (C_ipd(2)'last_event,  tpd_C_O((511 - 10)- 32*13 ), true),
						38 => (C_ipd(3)'last_event,  tpd_C_O((511 - 10)- 32*12 ), true),
						39=> (C_ipd(4)'last_event,  tpd_C_O((511 - 10)- 32*11 ), true), 
						40=> (C_ipd(5)'last_event,  tpd_C_O((511 - 10)- 32*10 ), true),
						41 => (C_ipd(6)'last_event,  tpd_C_O((511 - 10)- 32*9 ), true),
						42 => (C_ipd(7)'last_event,  tpd_C_O((511 - 10)- 32*8 ), true),
						43=> (C_ipd(8)'last_event,  tpd_C_O((511 - 10)- 32*7), true),
						44 => (C_ipd(9)'last_event,  tpd_C_O((511 - 10)- 32*6 ), true),
						45=> (C_ipd(10)'last_event,  tpd_C_O((511 - 10)- 32*5 ), true),
						46 => (C_ipd(11)'last_event,  tpd_C_O((511 - 10)- 32*4 ), true),
						47 => (C_ipd(12)'last_event,  tpd_C_O((511 - 10)- 32*3 ), true),
						48=> (C_ipd(13)'last_event,  tpd_C_O((511 - 10)- 32*2 ), true),
						49=> (C_ipd(14)'last_event,  tpd_C_O((511 - 10)- 32*1 ), true), 
						50=> (C_ipd(15)'last_event,  tpd_C_O((511 - 10)- 32*0 ), true),
						51=> (D_ipd(0)'last_event,  tpd_D_O((511 - 10)- 32*15 ), true),
						52 => (D_ipd(1)'last_event,  tpd_D_O((511 - 10)- 32*14 ), true),
						53 => (D_ipd(2)'last_event,  tpd_D_O((511 - 10)- 32*13 ), true),
						54 => (D_ipd(3)'last_event,  tpd_D_O((511 - 10)- 32*12 ), true),
						55=> (D_ipd(4)'last_event,  tpd_D_O((511 - 10)- 32*11 ), true), 
						56=> (D_ipd(5)'last_event,  tpd_D_O((511 - 10)- 32*10 ), true),
						57 => (D_ipd(6)'last_event,  tpd_D_O((511 - 10)- 32*9 ), true),
						58 => (D_ipd(7)'last_event,  tpd_D_O((511 - 10)- 32*8 ), true),
						59=> (D_ipd(8)'last_event,  tpd_D_O((511 - 10)- 32*7 ), true),
						60 => (D_ipd(9)'last_event,  tpd_D_O((511 - 10)- 32*6 ), true),
						61=> (D_ipd(10)'last_event,  tpd_D_O((511 - 10)- 32*5 ), true),
						62 => (D_ipd(11)'last_event,  tpd_D_O((511 - 10)- 32*4 ), true),
						63 => (D_ipd(12)'last_event,  tpd_D_O((511 - 10)- 32*3 ), true),
						64=> (D_ipd(13)'last_event,  tpd_D_O((511 - 10)- 32*2 ), true),
						65=> (D_ipd(14)'last_event,  tpd_D_O((511 - 10)- 32*1 ), true), 
						66=> (D_ipd(15)'last_event,  tpd_D_O((511 - 10)- 32*0 ), true),
						67=> (CI_ipd'last_event, tpd_CI_O(21), true)  ,  
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(21), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(21),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(21),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(21),true)),
      Mode          => VitalTransport,
	  IgnoreDefaultDelay => TRUE, 
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);   
	  
	  
	  	  	  	   VitalPathDelay01 (
      OutSignal     => O(22),
      GlitchData    => O_GlitchData(22),
      OutSignalName => "O(22)",
      OutTemp       => O_zd(22),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(22), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(22), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(22), true),
							3 => (A_ipd(0)'last_event,  tpd_A_O((511 - 9)- 32*15 ), true),
						4 => (A_ipd(1)'last_event,  tpd_A_O((511 - 9)- 32*14 ), true),
						5 => (A_ipd(2)'last_event,  tpd_A_O((511 - 9)- 32*13 ), true),
						6 => (A_ipd(3)'last_event,  tpd_A_O((511 - 9)- 32*12 ), true),
						7 => (A_ipd(4)'last_event,  tpd_A_O((511 - 9)- 32*11 ), true), 
						8 => (A_ipd(5)'last_event,  tpd_A_O((511 - 9)- 32*10 ), true),
						9 => (A_ipd(6)'last_event,  tpd_A_O((511 - 9)- 32*9 ), true),
						10 => (A_ipd(7)'last_event,  tpd_A_O((511 - 9)- 32*8 ), true),
						11=> (A_ipd(8)'last_event,  tpd_A_O((511 - 9)- 32*7 ), true),
						12 => (A_ipd(9)'last_event,  tpd_A_O((511 - 9)- 32*6 ), true),
						13 => (A_ipd(10)'last_event,  tpd_A_O((511 - 9)- 32*5 ), true),
						14 => (A_ipd(11)'last_event,  tpd_A_O((511 - 9)- 32*4 ), true),
						15 => (A_ipd(12)'last_event,  tpd_A_O((511 - 9)- 32*3 ), true),
						16=> (A_ipd(13)'last_event,  tpd_A_O((511 - 9)- 32*2), true),
						17=> (A_ipd(14)'last_event,  tpd_A_O((511 - 9)- 32*1 ), true), 
						18=> (A_ipd(15)'last_event,  tpd_A_O((511 - 9)- 32*0 ), true), 
						19=> (B_ipd(0)'last_event,  tpd_B_O((511 - 9)- 32*15 ), true),
						20 => (B_ipd(1)'last_event,  tpd_B_O((511 - 9)- 32*14 ), true),
						21 => (B_ipd(2)'last_event,  tpd_B_O((511 - 9)- 32*13 ), true),
						22 => (B_ipd(3)'last_event,  tpd_B_O((511 - 9)- 32*12 ), true),
						23=> (B_ipd(4)'last_event,  tpd_B_O((511 - 9)- 32*11 ), true), 
						24=> (B_ipd(5)'last_event,  tpd_B_O((511 - 9)- 32*10 ), true),
						25 => (B_ipd(6)'last_event,  tpd_B_O((511 - 9)- 32*9 ), true),
						26 => (B_ipd(7)'last_event,  tpd_B_O((511 - 9)- 32*8 ), true),
						27=> (B_ipd(8)'last_event,  tpd_B_O((511 - 9)- 32*7), true),
						28 => (B_ipd(9)'last_event,  tpd_B_O((511 - 9)- 32*6 ), true),
						29=> (B_ipd(10)'last_event,  tpd_B_O((511 - 9)- 32*5 ), true),
						30 => (B_ipd(11)'last_event,  tpd_B_O((511 - 9)- 32*4 ), true),
						31 => (B_ipd(12)'last_event,  tpd_B_O((511 - 9)- 32*3 ), true),
						32=> (B_ipd(13)'last_event,  tpd_B_O((511 - 9)- 32*2 ), true),
						33=> (B_ipd(14)'last_event,  tpd_B_O((511 - 9)- 32*1 ), true), 
						34=> (B_ipd(15)'last_event,  tpd_B_O((511 - 9)- 32*0 ), true),
						35=> (C_ipd(0)'last_event,  tpd_C_O((511 - 9)- 32*15 ), true),
						36 => (C_ipd(1)'last_event,  tpd_C_O((511 - 9)- 32*14 ), true),
						37 => (C_ipd(2)'last_event,  tpd_C_O((511 - 9)- 32*13 ), true),
						38 => (C_ipd(3)'last_event,  tpd_C_O((511 - 9)- 32*12 ), true),
						39=> (C_ipd(4)'last_event,  tpd_C_O((511 - 9)- 32*11 ), true), 
						40=> (C_ipd(5)'last_event,  tpd_C_O((511 - 9)- 32*10 ), true),
						41 => (C_ipd(6)'last_event,  tpd_C_O((511 - 9)- 32*9 ), true),
						42 => (C_ipd(7)'last_event,  tpd_C_O((511 - 9)- 32*8 ), true),
						43=> (C_ipd(8)'last_event,  tpd_C_O((511 - 9)- 32*7), true),
						44 => (C_ipd(9)'last_event,  tpd_C_O((511 - 9)- 32*6 ), true),
						45=> (C_ipd(10)'last_event,  tpd_C_O((511 - 9)- 32*5 ), true),
						46 => (C_ipd(11)'last_event,  tpd_C_O((511 - 9)- 32*4 ), true),
						47 => (C_ipd(12)'last_event,  tpd_C_O((511 - 9)- 32*3 ), true),
						48=> (C_ipd(13)'last_event,  tpd_C_O((511 - 9)- 32*2 ), true),
						49=> (C_ipd(14)'last_event,  tpd_C_O((511 - 9)- 32*1 ), true), 
						50=> (C_ipd(15)'last_event,  tpd_C_O((511 - 9)- 32*0 ), true),
						51=> (D_ipd(0)'last_event,  tpd_D_O((511 - 9)- 32*15 ), true),
						52 => (D_ipd(1)'last_event,  tpd_D_O((511 - 9)- 32*14 ), true),
						53 => (D_ipd(2)'last_event,  tpd_D_O((511 - 9)- 32*13 ), true),
						54 => (D_ipd(3)'last_event,  tpd_D_O((511 - 9)- 32*12 ), true),
						55=> (D_ipd(4)'last_event,  tpd_D_O((511 - 9)- 32*11 ), true), 
						56=> (D_ipd(5)'last_event,  tpd_D_O((511 - 9)- 32*10 ), true),
						57 => (D_ipd(6)'last_event,  tpd_D_O((511 - 9)- 32*9 ), true),
						58 => (D_ipd(7)'last_event,  tpd_D_O((511 - 9)- 32*8 ), true),
						59=> (D_ipd(8)'last_event,  tpd_D_O((511 - 9)- 32*7 ), true),
						60 => (D_ipd(9)'last_event,  tpd_D_O((511 - 9)- 32*6 ), true),
						61=> (D_ipd(10)'last_event,  tpd_D_O((511 - 9)- 32*5 ), true),
						62 => (D_ipd(11)'last_event,  tpd_D_O((511 - 9)- 32*4 ), true),
						63 => (D_ipd(12)'last_event,  tpd_D_O((511 - 9)- 32*3 ), true),
						64=> (D_ipd(13)'last_event,  tpd_D_O((511 - 9)- 32*2 ), true),
						65=> (D_ipd(14)'last_event,  tpd_D_O((511 - 9)- 32*1 ), true), 
						66=> (D_ipd(15)'last_event,  tpd_D_O((511 - 9)- 32*0 ), true),
						67=> (CI_ipd'last_event, tpd_CI_O(22), true)  ,  
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(22), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(22),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(22),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(22),true)),
      Mode          => VitalTransport,	  
	  IgnoreDefaultDelay => TRUE,		
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);  		
	  
	  
	  
	  	  	  	   VitalPathDelay01 (
      OutSignal     => O(23),
      GlitchData    => O_GlitchData(23),
      OutSignalName => "O(23)",
      OutTemp       => O_zd(23),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(23), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(23), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(23), true),
							3 => (A_ipd(0)'last_event,  tpd_A_O((511 - 8)- 32*15 ), true),
						4 => (A_ipd(1)'last_event,  tpd_A_O((511 - 8)- 32*14 ), true),
						5 => (A_ipd(2)'last_event,  tpd_A_O((511 - 8)- 32*13 ), true),
						6 => (A_ipd(3)'last_event,  tpd_A_O((511 - 8)- 32*12 ), true),
						7 => (A_ipd(4)'last_event,  tpd_A_O((511 - 8)- 32*11 ), true), 
						8 => (A_ipd(5)'last_event,  tpd_A_O((511 - 8)- 32*10 ), true),
						9 => (A_ipd(6)'last_event,  tpd_A_O((511 - 8)- 32*9 ), true),
						10 => (A_ipd(7)'last_event,  tpd_A_O((511 - 8)- 32*8 ), true),
						11=> (A_ipd(8)'last_event,  tpd_A_O((511 - 8)- 32*7 ), true),
						12 => (A_ipd(9)'last_event,  tpd_A_O((511 - 8)- 32*6 ), true),
						13 => (A_ipd(10)'last_event,  tpd_A_O((511 - 8)- 32*5 ), true),
						14 => (A_ipd(11)'last_event,  tpd_A_O((511 - 8)- 32*4 ), true),
						15 => (A_ipd(12)'last_event,  tpd_A_O((511 - 8)- 32*3 ), true),
						16=> (A_ipd(13)'last_event,  tpd_A_O((511 - 8)- 32*2), true),
						17=> (A_ipd(14)'last_event,  tpd_A_O((511 - 8)- 32*1 ), true), 
						18=> (A_ipd(15)'last_event,  tpd_A_O((511 - 8)- 32*0 ), true), 
						19=> (B_ipd(0)'last_event,  tpd_B_O((511 - 8)- 32*15 ), true),
						20 => (B_ipd(1)'last_event,  tpd_B_O((511 - 8)- 32*14 ), true),
						21 => (B_ipd(2)'last_event,  tpd_B_O((511 - 8)- 32*13 ), true),
						22 => (B_ipd(3)'last_event,  tpd_B_O((511 - 8)- 32*12 ), true),
						23=> (B_ipd(4)'last_event,  tpd_B_O((511 - 8)- 32*11 ), true), 
						24=> (B_ipd(5)'last_event,  tpd_B_O((511 - 8)- 32*10 ), true),
						25 => (B_ipd(6)'last_event,  tpd_B_O((511 - 8)- 32*9 ), true),
						26 => (B_ipd(7)'last_event,  tpd_B_O((511 - 8)- 32*8 ), true),
						27=> (B_ipd(8)'last_event,  tpd_B_O((511 - 8)- 32*7), true),
						28 => (B_ipd(9)'last_event,  tpd_B_O((511 - 8)- 32*6 ), true),
						29=> (B_ipd(10)'last_event,  tpd_B_O((511 - 8)- 32*5 ), true),
						30 => (B_ipd(11)'last_event,  tpd_B_O((511 - 8)- 32*4 ), true),
						31 => (B_ipd(12)'last_event,  tpd_B_O((511 - 8)- 32*3 ), true),
						32=> (B_ipd(13)'last_event,  tpd_B_O((511 - 8)- 32*2 ), true),
						33=> (B_ipd(14)'last_event,  tpd_B_O((511 - 8)- 32*1 ), true), 
						34=> (B_ipd(15)'last_event,  tpd_B_O((511 - 8)- 32*0 ), true),
						35=> (C_ipd(0)'last_event,  tpd_C_O((511 - 8)- 32*15 ), true),
						36 => (C_ipd(1)'last_event,  tpd_C_O((511 - 8)- 32*14 ), true),
						37 => (C_ipd(2)'last_event,  tpd_C_O((511 - 8)- 32*13 ), true),
						38 => (C_ipd(3)'last_event,  tpd_C_O((511 - 8)- 32*12 ), true),
						39=> (C_ipd(4)'last_event,  tpd_C_O((511 - 8)- 32*11 ), true), 
						40=> (C_ipd(5)'last_event,  tpd_C_O((511 - 8)- 32*10 ), true),
						41 => (C_ipd(6)'last_event,  tpd_C_O((511 - 8)- 32*9 ), true),
						42 => (C_ipd(7)'last_event,  tpd_C_O((511 - 8)- 32*8 ), true),
						43=> (C_ipd(8)'last_event,  tpd_C_O((511 - 8)- 32*7), true),
						44 => (C_ipd(9)'last_event,  tpd_C_O((511 - 8)- 32*6 ), true),
						45=> (C_ipd(10)'last_event,  tpd_C_O((511 - 8)- 32*5 ), true),
						46 => (C_ipd(11)'last_event,  tpd_C_O((511 - 8)- 32*4 ), true),
						47 => (C_ipd(12)'last_event,  tpd_C_O((511 - 8)- 32*3 ), true),
						48=> (C_ipd(13)'last_event,  tpd_C_O((511 - 8)- 32*2 ), true),
						49=> (C_ipd(14)'last_event,  tpd_C_O((511 - 8)- 32*1 ), true), 
						50=> (C_ipd(15)'last_event,  tpd_C_O((511 - 8)- 32*0 ), true),
						51=> (D_ipd(0)'last_event,  tpd_D_O((511 - 8)- 32*15 ), true),
						52 => (D_ipd(1)'last_event,  tpd_D_O((511 - 8)- 32*14 ), true),
						53 => (D_ipd(2)'last_event,  tpd_D_O((511 - 8)- 32*13 ), true),
						54 => (D_ipd(3)'last_event,  tpd_D_O((511 - 8)- 32*12 ), true),
						55=> (D_ipd(4)'last_event,  tpd_D_O((511 - 8)- 32*11 ), true), 
						56=> (D_ipd(5)'last_event,  tpd_D_O((511 - 8)- 32*10 ), true),
						57 => (D_ipd(6)'last_event,  tpd_D_O((511 - 8)- 32*9 ), true),
						58 => (D_ipd(7)'last_event,  tpd_D_O((511 - 8)- 32*8 ), true),
						59=> (D_ipd(8)'last_event,  tpd_D_O((511 - 8)- 32*7 ), true),
						60 => (D_ipd(9)'last_event,  tpd_D_O((511 - 8)- 32*6 ), true),
						61=> (D_ipd(10)'last_event,  tpd_D_O((511 - 8)- 32*5 ), true),
						62 => (D_ipd(11)'last_event,  tpd_D_O((511 - 8)- 32*4 ), true),
						63 => (D_ipd(12)'last_event,  tpd_D_O((511 - 8)- 32*3 ), true),
						64=> (D_ipd(13)'last_event,  tpd_D_O((511 - 8)- 32*2 ), true),
						65=> (D_ipd(14)'last_event,  tpd_D_O((511 - 8)- 32*1 ), true), 
						66=> (D_ipd(15)'last_event,  tpd_D_O((511 - 8)- 32*0 ), true),
						67=> (CI_ipd'last_event, tpd_CI_O(23), true)  ,  
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(23), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(23),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(23),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(23),true)),
      Mode          => VitalTransport,	   
	  IgnoreDefaultDelay => TRUE,
      RejectFastPath=>TRUE,
	  Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);  		
	  
	  
	  
	  	  	  	   VitalPathDelay01 (
      OutSignal     => O(24),
      GlitchData    => O_GlitchData(24),
      OutSignalName => "O(24)",
      OutTemp       => O_zd(24),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(24), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(24), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(24), true),
						3 => (A_ipd(0)'last_event,  tpd_A_O((511 - 7)- 32*15 ), true),
						4 => (A_ipd(1)'last_event,  tpd_A_O((511 - 7)- 32*14 ), true),
						5 => (A_ipd(2)'last_event,  tpd_A_O((511 - 7)- 32*13 ), true),
						6 => (A_ipd(3)'last_event,  tpd_A_O((511 - 7)- 32*12 ), true),
						7 => (A_ipd(4)'last_event,  tpd_A_O((511 - 7)- 32*11 ), true), 
						8 => (A_ipd(5)'last_event,  tpd_A_O((511 - 7)- 32*10 ), true),
						9 => (A_ipd(6)'last_event,  tpd_A_O((511 - 7)- 32*9 ), true),
						10 => (A_ipd(7)'last_event,  tpd_A_O((511 - 7)- 32*8 ), true),
						11=> (A_ipd(8)'last_event,  tpd_A_O((511 - 7)- 32*7 ), true),
						12 => (A_ipd(9)'last_event,  tpd_A_O((511 - 7)- 32*6 ), true),
						13 => (A_ipd(10)'last_event,  tpd_A_O((511 - 7)- 32*5 ), true),
						14 => (A_ipd(11)'last_event,  tpd_A_O((511 - 7)- 32*4 ), true),
						15 => (A_ipd(12)'last_event,  tpd_A_O((511 - 7)- 32*3 ), true),
						16=> (A_ipd(13)'last_event,  tpd_A_O((511 - 7)- 32*2), true),
						17=> (A_ipd(14)'last_event,  tpd_A_O((511 - 7)- 32*1 ), true), 
						18=> (A_ipd(15)'last_event,  tpd_A_O((511 - 7)- 32*0 ), true), 
						19=> (B_ipd(0)'last_event,  tpd_B_O((511 - 7)- 32*15 ), true),
						20 => (B_ipd(1)'last_event,  tpd_B_O((511 - 7)- 32*14 ), true),
						21 => (B_ipd(2)'last_event,  tpd_B_O((511 - 7)- 32*13 ), true),
						22 => (B_ipd(3)'last_event,  tpd_B_O((511 - 7)- 32*12 ), true),
						23=> (B_ipd(4)'last_event,  tpd_B_O((511 - 7)- 32*11 ), true), 
						24=> (B_ipd(5)'last_event,  tpd_B_O((511 - 7)- 32*10 ), true),
						25 => (B_ipd(6)'last_event,  tpd_B_O((511 - 7)- 32*9 ), true),
						26 => (B_ipd(7)'last_event,  tpd_B_O((511 - 7)- 32*8 ), true),
						27=> (B_ipd(8)'last_event,  tpd_B_O((511 - 7)- 32*7), true),
						28 => (B_ipd(9)'last_event,  tpd_B_O((511 - 7)- 32*6 ), true),
						29=> (B_ipd(10)'last_event,  tpd_B_O((511 - 7)- 32*5 ), true),
						30 => (B_ipd(11)'last_event,  tpd_B_O((511 - 7)- 32*4 ), true),
						31 => (B_ipd(12)'last_event,  tpd_B_O((511 - 7)- 32*3 ), true),
						32=> (B_ipd(13)'last_event,  tpd_B_O((511 - 7)- 32*2 ), true),
						33=> (B_ipd(14)'last_event,  tpd_B_O((511 - 7)- 32*1 ), true), 
						34=> (B_ipd(15)'last_event,  tpd_B_O((511 - 7)- 32*0 ), true),
						35=> (C_ipd(0)'last_event,  tpd_C_O((511 - 7)- 32*15 ), true),
						36 => (C_ipd(1)'last_event,  tpd_C_O((511 - 7)- 32*14 ), true),
						37 => (C_ipd(2)'last_event,  tpd_C_O((511 - 7)- 32*13 ), true),
						38 => (C_ipd(3)'last_event,  tpd_C_O((511 - 7)- 32*12 ), true),
						39=> (C_ipd(4)'last_event,  tpd_C_O((511 - 7)- 32*11 ), true), 
						40=> (C_ipd(5)'last_event,  tpd_C_O((511 - 7)- 32*10 ), true),
						41 => (C_ipd(6)'last_event,  tpd_C_O((511 - 7)- 32*9 ), true),
						42 => (C_ipd(7)'last_event,  tpd_C_O((511 - 7)- 32*8 ), true),
						43=> (C_ipd(8)'last_event,  tpd_C_O((511 - 7)- 32*7), true),
						44 => (C_ipd(9)'last_event,  tpd_C_O((511 - 7)- 32*6 ), true),
						45=> (C_ipd(10)'last_event,  tpd_C_O((511 - 7)- 32*5 ), true),
						46 => (C_ipd(11)'last_event,  tpd_C_O((511 - 7)- 32*4 ), true),
						47 => (C_ipd(12)'last_event,  tpd_C_O((511 - 7)- 32*3 ), true),
						48=> (C_ipd(13)'last_event,  tpd_C_O((511 - 7)- 32*2 ), true),
						49=> (C_ipd(14)'last_event,  tpd_C_O((511 - 7)- 32*1 ), true), 
						50=> (C_ipd(15)'last_event,  tpd_C_O((511 - 7)- 32*0 ), true),
						51=> (D_ipd(0)'last_event,  tpd_D_O((511 - 7)- 32*15 ), true),
						52 => (D_ipd(1)'last_event,  tpd_D_O((511 - 7)- 32*14 ), true),
						53 => (D_ipd(2)'last_event,  tpd_D_O((511 - 7)- 32*13 ), true),
						54 => (D_ipd(3)'last_event,  tpd_D_O((511 - 7)- 32*12 ), true),
						55=> (D_ipd(4)'last_event,  tpd_D_O((511 - 7)- 32*11 ), true), 
						56=> (D_ipd(5)'last_event,  tpd_D_O((511 - 7)- 32*10 ), true),
						57 => (D_ipd(6)'last_event,  tpd_D_O((511 - 7)- 32*9 ), true),
						58 => (D_ipd(7)'last_event,  tpd_D_O((511 - 7)- 32*8 ), true),
						59=> (D_ipd(8)'last_event,  tpd_D_O((511 - 7)- 32*7 ), true),
						60 => (D_ipd(9)'last_event,  tpd_D_O((511 - 7)- 32*6 ), true),
						61=> (D_ipd(10)'last_event,  tpd_D_O((511 - 7)- 32*5 ), true),
						62 => (D_ipd(11)'last_event,  tpd_D_O((511 - 7)- 32*4 ), true),
						63 => (D_ipd(12)'last_event,  tpd_D_O((511 - 7)- 32*3 ), true),
						64=> (D_ipd(13)'last_event,  tpd_D_O((511 - 7)- 32*2 ), true),
						65=> (D_ipd(14)'last_event,  tpd_D_O((511 - 7)- 32*1 ), true), 
						66=> (D_ipd(15)'last_event,  tpd_D_O((511 - 7)- 32*0 ), true),
						67=> (CI_ipd'last_event, tpd_CI_O(24), true)  ,  
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(24), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(24),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(24),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(24),true)),
      Mode          => VitalTransport,	
	  IgnoreDefaultDelay => TRUE,	  
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);  
	  
	  
	  
	  	  	  	   VitalPathDelay01 (
      OutSignal     => O(25),
      GlitchData    => O_GlitchData(25),
      OutSignalName => "O(25)",
      OutTemp       => O_zd(25),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(25), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(25), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(25), true),
							3 => (A_ipd(0)'last_event,  tpd_A_O((511 - 6)- 32*15 ), true),
						4 => (A_ipd(1)'last_event,  tpd_A_O((511 - 6)- 32*14 ), true),
						5 => (A_ipd(2)'last_event,  tpd_A_O((511 - 6)- 32*13 ), true),
						6 => (A_ipd(3)'last_event,  tpd_A_O((511 - 6)- 32*12 ), true),
						7 => (A_ipd(4)'last_event,  tpd_A_O((511 - 6)- 32*11 ), true), 
						8 => (A_ipd(5)'last_event,  tpd_A_O((511 - 6)- 32*10 ), true),
						9 => (A_ipd(6)'last_event,  tpd_A_O((511 - 6)- 32*9 ), true),
						10 => (A_ipd(7)'last_event,  tpd_A_O((511 - 6)- 32*8 ), true),
						11=> (A_ipd(8)'last_event,  tpd_A_O((511 - 6)- 32*7 ), true),
						12 => (A_ipd(9)'last_event,  tpd_A_O((511 - 6)- 32*6 ), true),
						13 => (A_ipd(10)'last_event,  tpd_A_O((511 - 6)- 32*5 ), true),
						14 => (A_ipd(11)'last_event,  tpd_A_O((511 - 6)- 32*4 ), true),
						15 => (A_ipd(12)'last_event,  tpd_A_O((511 - 6)- 32*3 ), true),
						16=> (A_ipd(13)'last_event,  tpd_A_O((511 - 6)- 32*2), true),
						17=> (A_ipd(14)'last_event,  tpd_A_O((511 - 6)- 32*1 ), true), 
						18=> (A_ipd(15)'last_event,  tpd_A_O((511 - 6)- 32*0 ), true), 
						19=> (B_ipd(0)'last_event,  tpd_B_O((511 - 6)- 32*15 ), true),
						20 => (B_ipd(1)'last_event,  tpd_B_O((511 - 6)- 32*14 ), true),
						21 => (B_ipd(2)'last_event,  tpd_B_O((511 - 6)- 32*13 ), true),
						22 => (B_ipd(3)'last_event,  tpd_B_O((511 - 6)- 32*12 ), true),
						23=> (B_ipd(4)'last_event,  tpd_B_O((511 - 6)- 32*11 ), true), 
						24=> (B_ipd(5)'last_event,  tpd_B_O((511 - 6)- 32*10 ), true),
						25 => (B_ipd(6)'last_event,  tpd_B_O((511 - 6)- 32*9 ), true),
						26 => (B_ipd(7)'last_event,  tpd_B_O((511 - 6)- 32*8 ), true),
						27=> (B_ipd(8)'last_event,  tpd_B_O((511 - 6)- 32*7), true),
						28 => (B_ipd(9)'last_event,  tpd_B_O((511 - 6)- 32*6 ), true),
						29=> (B_ipd(10)'last_event,  tpd_B_O((511 - 6)- 32*5 ), true),
						30 => (B_ipd(11)'last_event,  tpd_B_O((511 - 6)- 32*4 ), true),
						31 => (B_ipd(12)'last_event,  tpd_B_O((511 - 6)- 32*3 ), true),
						32=> (B_ipd(13)'last_event,  tpd_B_O((511 - 6)- 32*2 ), true),
						33=> (B_ipd(14)'last_event,  tpd_B_O((511 - 6)- 32*1 ), true), 
						34=> (B_ipd(15)'last_event,  tpd_B_O((511 - 6)- 32*0 ), true),
						35=> (C_ipd(0)'last_event,  tpd_C_O((511 - 6)- 32*15 ), true),
						36 => (C_ipd(1)'last_event,  tpd_C_O((511 - 6)- 32*14 ), true),
						37 => (C_ipd(2)'last_event,  tpd_C_O((511 - 6)- 32*13 ), true),
						38 => (C_ipd(3)'last_event,  tpd_C_O((511 - 6)- 32*12 ), true),
						39=> (C_ipd(4)'last_event,  tpd_C_O((511 - 6)- 32*11 ), true), 
						40=> (C_ipd(5)'last_event,  tpd_C_O((511 - 6)- 32*10 ), true),
						41 => (C_ipd(6)'last_event,  tpd_C_O((511 - 6)- 32*9 ), true),
						42 => (C_ipd(7)'last_event,  tpd_C_O((511 - 6)- 32*8 ), true),
						43=> (C_ipd(8)'last_event,  tpd_C_O((511 - 6)- 32*7), true),
						44 => (C_ipd(9)'last_event,  tpd_C_O((511 - 6)- 32*6 ), true),
						45=> (C_ipd(10)'last_event,  tpd_C_O((511 - 6)- 32*5 ), true),
						46 => (C_ipd(11)'last_event,  tpd_C_O((511 - 6)- 32*4 ), true),
						47 => (C_ipd(12)'last_event,  tpd_C_O((511 - 6)- 32*3 ), true),
						48=> (C_ipd(13)'last_event,  tpd_C_O((511 - 6)- 32*2 ), true),
						49=> (C_ipd(14)'last_event,  tpd_C_O((511 - 6)- 32*1 ), true), 
						50=> (C_ipd(15)'last_event,  tpd_C_O((511 - 6)- 32*0 ), true),
						51=> (D_ipd(0)'last_event,  tpd_D_O((511 - 6)- 32*15 ), true),
						52 => (D_ipd(1)'last_event,  tpd_D_O((511 - 6)- 32*14 ), true),
						53 => (D_ipd(2)'last_event,  tpd_D_O((511 - 6)- 32*13 ), true),
						54 => (D_ipd(3)'last_event,  tpd_D_O((511 - 6)- 32*12 ), true),
						55=> (D_ipd(4)'last_event,  tpd_D_O((511 - 6)- 32*11 ), true), 
						56=> (D_ipd(5)'last_event,  tpd_D_O((511 - 6)- 32*10 ), true),
						57 => (D_ipd(6)'last_event,  tpd_D_O((511 - 6)- 32*9 ), true),
						58 => (D_ipd(7)'last_event,  tpd_D_O((511 - 6)- 32*8 ), true),
						59=> (D_ipd(8)'last_event,  tpd_D_O((511 - 6)- 32*7 ), true),
						60 => (D_ipd(9)'last_event,  tpd_D_O((511 - 6)- 32*6 ), true),
						61=> (D_ipd(10)'last_event,  tpd_D_O((511 - 6)- 32*5 ), true),
						62 => (D_ipd(11)'last_event,  tpd_D_O((511 - 6)- 32*4 ), true),
						63 => (D_ipd(12)'last_event,  tpd_D_O((511 - 6)- 32*3 ), true),
						64=> (D_ipd(13)'last_event,  tpd_D_O((511 - 6)- 32*2 ), true),
						65=> (D_ipd(14)'last_event,  tpd_D_O((511 - 6)- 32*1 ), true), 
						66=> (D_ipd(15)'last_event,  tpd_D_O((511 - 6)- 32*0 ), true),
						67=> (CI_ipd'last_event, tpd_CI_O(25), true)  ,  
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(25), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(25),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(25),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(25),true)),
      Mode          => VitalTransport,
	  IgnoreDefaultDelay => TRUE,	   
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);  
	  
	  
	  
	  
	  	  	  	   VitalPathDelay01 (
      OutSignal     => O(26),
      GlitchData    => O_GlitchData(26),
      OutSignalName => "O(26)",
      OutTemp       => O_zd(26),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(26), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(26), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(26), true),
							3 => (A_ipd(0)'last_event,  tpd_A_O((511 - 5)- 32*15 ), true),
						4 => (A_ipd(1)'last_event,  tpd_A_O((511 - 5)- 32*14 ), true),
						5 => (A_ipd(2)'last_event,  tpd_A_O((511 - 5)- 32*13 ), true),
						6 => (A_ipd(3)'last_event,  tpd_A_O((511 - 5)- 32*12 ), true),
						7 => (A_ipd(4)'last_event,  tpd_A_O((511 - 5)- 32*11 ), true), 
						8 => (A_ipd(5)'last_event,  tpd_A_O((511 - 5)- 32*10 ), true),
						9 => (A_ipd(6)'last_event,  tpd_A_O((511 - 5)- 32*9 ), true),
						10 => (A_ipd(7)'last_event,  tpd_A_O((511 - 5)- 32*8 ), true),
						11=> (A_ipd(8)'last_event,  tpd_A_O((511 - 5)- 32*7 ), true),
						12 => (A_ipd(9)'last_event,  tpd_A_O((511 - 5)- 32*6 ), true),
						13 => (A_ipd(10)'last_event,  tpd_A_O((511 - 5)- 32*5 ), true),
						14 => (A_ipd(11)'last_event,  tpd_A_O((511 - 5)- 32*4 ), true),
						15 => (A_ipd(12)'last_event,  tpd_A_O((511 - 5)- 32*3 ), true),
						16=> (A_ipd(13)'last_event,  tpd_A_O((511 - 5)- 32*2), true),
						17=> (A_ipd(14)'last_event,  tpd_A_O((511 - 5)- 32*1 ), true), 
						18=> (A_ipd(15)'last_event,  tpd_A_O((511 - 5)- 32*0 ), true), 
						19=> (B_ipd(0)'last_event,  tpd_B_O((511 - 5)- 32*15 ), true),
						20 => (B_ipd(1)'last_event,  tpd_B_O((511 - 5)- 32*14 ), true),
						21 => (B_ipd(2)'last_event,  tpd_B_O((511 - 5)- 32*13 ), true),
						22 => (B_ipd(3)'last_event,  tpd_B_O((511 - 5)- 32*12 ), true),
						23=> (B_ipd(4)'last_event,  tpd_B_O((511 - 5)- 32*11 ), true), 
						24=> (B_ipd(5)'last_event,  tpd_B_O((511 - 5)- 32*10 ), true),
						25 => (B_ipd(6)'last_event,  tpd_B_O((511 - 5)- 32*9 ), true),
						26 => (B_ipd(7)'last_event,  tpd_B_O((511 - 5)- 32*8 ), true),
						27=> (B_ipd(8)'last_event,  tpd_B_O((511 - 5)- 32*7), true),
						28 => (B_ipd(9)'last_event,  tpd_B_O((511 - 5)- 32*6 ), true),
						29=> (B_ipd(10)'last_event,  tpd_B_O((511 - 5)- 32*5 ), true),
						30 => (B_ipd(11)'last_event,  tpd_B_O((511 - 5)- 32*4 ), true),
						31 => (B_ipd(12)'last_event,  tpd_B_O((511 - 5)- 32*3 ), true),
						32=> (B_ipd(13)'last_event,  tpd_B_O((511 - 5)- 32*2 ), true),
						33=> (B_ipd(14)'last_event,  tpd_B_O((511 - 5)- 32*1 ), true), 
						34=> (B_ipd(15)'last_event,  tpd_B_O((511 - 5)- 32*0 ), true),
						35=> (C_ipd(0)'last_event,  tpd_C_O((511 - 5)- 32*15 ), true),
						36 => (C_ipd(1)'last_event,  tpd_C_O((511 - 5)- 32*14 ), true),
						37 => (C_ipd(2)'last_event,  tpd_C_O((511 - 5)- 32*13 ), true),
						38 => (C_ipd(3)'last_event,  tpd_C_O((511 - 5)- 32*12 ), true),
						39=> (C_ipd(4)'last_event,  tpd_C_O((511 - 5)- 32*11 ), true), 
						40=> (C_ipd(5)'last_event,  tpd_C_O((511 - 5)- 32*10 ), true),
						41 => (C_ipd(6)'last_event,  tpd_C_O((511 - 5)- 32*9 ), true),
						42 => (C_ipd(7)'last_event,  tpd_C_O((511 - 5)- 32*8 ), true),
						43=> (C_ipd(8)'last_event,  tpd_C_O((511 - 5)- 32*7), true),
						44 => (C_ipd(9)'last_event,  tpd_C_O((511 - 5)- 32*6 ), true),
						45=> (C_ipd(10)'last_event,  tpd_C_O((511 - 5)- 32*5 ), true),
						46 => (C_ipd(11)'last_event,  tpd_C_O((511 - 5)- 32*4 ), true),
						47 => (C_ipd(12)'last_event,  tpd_C_O((511 - 5)- 32*3 ), true),
						48=> (C_ipd(13)'last_event,  tpd_C_O((511 - 5)- 32*2 ), true),
						49=> (C_ipd(14)'last_event,  tpd_C_O((511 - 5)- 32*1 ), true), 
						50=> (C_ipd(15)'last_event,  tpd_C_O((511 - 5)- 32*0 ), true),
						51=> (D_ipd(0)'last_event,  tpd_D_O((511 - 5)- 32*15 ), true),
						52 => (D_ipd(1)'last_event,  tpd_D_O((511 - 5)- 32*14 ), true),
						53 => (D_ipd(2)'last_event,  tpd_D_O((511 - 5)- 32*13 ), true),
						54 => (D_ipd(3)'last_event,  tpd_D_O((511 - 5)- 32*12 ), true),
						55=> (D_ipd(4)'last_event,  tpd_D_O((511 - 5)- 32*11 ), true), 
						56=> (D_ipd(5)'last_event,  tpd_D_O((511 - 5)- 32*10 ), true),
						57 => (D_ipd(6)'last_event,  tpd_D_O((511 - 5)- 32*9 ), true),
						58 => (D_ipd(7)'last_event,  tpd_D_O((511 - 5)- 32*8 ), true),
						59=> (D_ipd(8)'last_event,  tpd_D_O((511 - 5)- 32*7 ), true),
						60 => (D_ipd(9)'last_event,  tpd_D_O((511 - 5)- 32*6 ), true),
						61=> (D_ipd(10)'last_event,  tpd_D_O((511 - 5)- 32*5 ), true),
						62 => (D_ipd(11)'last_event,  tpd_D_O((511 - 5)- 32*4 ), true),
						63 => (D_ipd(12)'last_event,  tpd_D_O((511 - 5)- 32*3 ), true),
						64=> (D_ipd(13)'last_event,  tpd_D_O((511 - 5)- 32*2 ), true),
						65=> (D_ipd(14)'last_event,  tpd_D_O((511 - 5)- 32*1 ), true), 
						66=> (D_ipd(15)'last_event,  tpd_D_O((511 - 5)- 32*0 ), true),
						67=> (CI_ipd'last_event, tpd_CI_O(26), true)  ,  
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(26), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(26),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(26),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(26),true)),
      Mode          => VitalTransport,		  
	  IgnoreDefaultDelay => TRUE,	  
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);  
	  
	  
	  
	  	  	  	   VitalPathDelay01 (
      OutSignal     => O(27),
      GlitchData    => O_GlitchData(27),
      OutSignalName => "O(27)",
      OutTemp       => O_zd(27),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(27), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(27), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(27), true),
							3 => (A_ipd(0)'last_event,  tpd_A_O((511 - 4)- 32*15 ), true),
						4 => (A_ipd(1)'last_event,  tpd_A_O((511 - 4)- 32*14 ), true),
						5 => (A_ipd(2)'last_event,  tpd_A_O((511 - 4)- 32*13 ), true),
						6 => (A_ipd(3)'last_event,  tpd_A_O((511 - 4)- 32*12 ), true),
						7 => (A_ipd(4)'last_event,  tpd_A_O((511 - 4)- 32*11 ), true), 
						8 => (A_ipd(5)'last_event,  tpd_A_O((511 - 4)- 32*10 ), true),
						9 => (A_ipd(6)'last_event,  tpd_A_O((511 - 4)- 32*9 ), true),
						10 => (A_ipd(7)'last_event,  tpd_A_O((511 - 4)- 32*8 ), true),
						11=> (A_ipd(8)'last_event,  tpd_A_O((511 - 4)- 32*7 ), true),
						12 => (A_ipd(9)'last_event,  tpd_A_O((511 - 4)- 32*6 ), true),
						13 => (A_ipd(10)'last_event,  tpd_A_O((511 - 4)- 32*5 ), true),
						14 => (A_ipd(11)'last_event,  tpd_A_O((511 - 4)- 32*4 ), true),
						15 => (A_ipd(12)'last_event,  tpd_A_O((511 - 4)- 32*3 ), true),
						16=> (A_ipd(13)'last_event,  tpd_A_O((511 - 4)- 32*2), true),
						17=> (A_ipd(14)'last_event,  tpd_A_O((511 - 4)- 32*1 ), true), 
						18=> (A_ipd(15)'last_event,  tpd_A_O((511 - 4)- 32*0 ), true), 
						19=> (B_ipd(0)'last_event,  tpd_B_O((511 - 4)- 32*15 ), true),
						20 => (B_ipd(1)'last_event,  tpd_B_O((511 - 4)- 32*14 ), true),
						21 => (B_ipd(2)'last_event,  tpd_B_O((511 - 4)- 32*13 ), true),
						22 => (B_ipd(3)'last_event,  tpd_B_O((511 - 4)- 32*12 ), true),
						23=> (B_ipd(4)'last_event,  tpd_B_O((511 - 4)- 32*11 ), true), 
						24=> (B_ipd(5)'last_event,  tpd_B_O((511 - 4)- 32*10 ), true),
						25 => (B_ipd(6)'last_event,  tpd_B_O((511 - 4)- 32*9 ), true),
						26 => (B_ipd(7)'last_event,  tpd_B_O((511 - 4)- 32*8 ), true),
						27=> (B_ipd(8)'last_event,  tpd_B_O((511 - 4)- 32*7), true),
						28 => (B_ipd(9)'last_event,  tpd_B_O((511 - 4)- 32*6 ), true),
						29=> (B_ipd(10)'last_event,  tpd_B_O((511 - 4)- 32*5 ), true),
						30 => (B_ipd(11)'last_event,  tpd_B_O((511 - 4)- 32*4 ), true),
						31 => (B_ipd(12)'last_event,  tpd_B_O((511 - 4)- 32*3 ), true),
						32=> (B_ipd(13)'last_event,  tpd_B_O((511 - 4)- 32*2 ), true),
						33=> (B_ipd(14)'last_event,  tpd_B_O((511 - 4)- 32*1 ), true), 
						34=> (B_ipd(15)'last_event,  tpd_B_O((511 - 4)- 32*0 ), true),
						35=> (C_ipd(0)'last_event,  tpd_C_O((511 - 4)- 32*15 ), true),
						36 => (C_ipd(1)'last_event,  tpd_C_O((511 - 4)- 32*14 ), true),
						37 => (C_ipd(2)'last_event,  tpd_C_O((511 - 4)- 32*13 ), true),
						38 => (C_ipd(3)'last_event,  tpd_C_O((511 - 4)- 32*12 ), true),
						39=> (C_ipd(4)'last_event,  tpd_C_O((511 - 4)- 32*11 ), true), 
						40=> (C_ipd(5)'last_event,  tpd_C_O((511 - 4)- 32*10 ), true),
						41 => (C_ipd(6)'last_event,  tpd_C_O((511 - 4)- 32*9 ), true),
						42 => (C_ipd(7)'last_event,  tpd_C_O((511 - 4)- 32*8 ), true),
						43=> (C_ipd(8)'last_event,  tpd_C_O((511 - 4)- 32*7), true),
						44 => (C_ipd(9)'last_event,  tpd_C_O((511 - 4)- 32*6 ), true),
						45=> (C_ipd(10)'last_event,  tpd_C_O((511 - 4)- 32*5 ), true),
						46 => (C_ipd(11)'last_event,  tpd_C_O((511 - 4)- 32*4 ), true),
						47 => (C_ipd(12)'last_event,  tpd_C_O((511 - 4)- 32*3 ), true),
						48=> (C_ipd(13)'last_event,  tpd_C_O((511 - 4)- 32*2 ), true),
						49=> (C_ipd(14)'last_event,  tpd_C_O((511 - 4)- 32*1 ), true), 
						50=> (C_ipd(15)'last_event,  tpd_C_O((511 - 4)- 32*0 ), true),
						51=> (D_ipd(0)'last_event,  tpd_D_O((511 - 4)- 32*15 ), true),
						52 => (D_ipd(1)'last_event,  tpd_D_O((511 - 4)- 32*14 ), true),
						53 => (D_ipd(2)'last_event,  tpd_D_O((511 - 4)- 32*13 ), true),
						54 => (D_ipd(3)'last_event,  tpd_D_O((511 - 4)- 32*12 ), true),
						55=> (D_ipd(4)'last_event,  tpd_D_O((511 - 4)- 32*11 ), true), 
						56=> (D_ipd(5)'last_event,  tpd_D_O((511 - 4)- 32*10 ), true),
						57 => (D_ipd(6)'last_event,  tpd_D_O((511 - 4)- 32*9 ), true),
						58 => (D_ipd(7)'last_event,  tpd_D_O((511 - 4)- 32*8 ), true),
						59=> (D_ipd(8)'last_event,  tpd_D_O((511 - 4)- 32*7 ), true),
						60 => (D_ipd(9)'last_event,  tpd_D_O((511 - 4)- 32*6 ), true),
						61=> (D_ipd(10)'last_event,  tpd_D_O((511 - 4)- 32*5 ), true),
						62 => (D_ipd(11)'last_event,  tpd_D_O((511 - 4)- 32*4 ), true),
						63 => (D_ipd(12)'last_event,  tpd_D_O((511 - 4)- 32*3 ), true),
						64=> (D_ipd(13)'last_event,  tpd_D_O((511 - 4)- 32*2 ), true),
						65=> (D_ipd(14)'last_event,  tpd_D_O((511 - 4)- 32*1 ), true), 
						66=> (D_ipd(15)'last_event,  tpd_D_O((511 - 4)- 32*0 ), true),
						67=> (CI_ipd'last_event, tpd_CI_O(27), true)  ,  
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(27), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(27),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(27),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(27),true)),
      Mode          => VitalTransport,		   
	  IgnoreDefaultDelay => TRUE,		 
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);  
	  
	  
	  
	  	  	  	   VitalPathDelay01 (
      OutSignal     => O(28),
      GlitchData    => O_GlitchData(28),
      OutSignalName => "O(28)",
      OutTemp       => O_zd(28),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(28), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(28), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(28), true),
							3 => (A_ipd(0)'last_event,  tpd_A_O((511 - 3)- 32*15 ), true),
						4 => (A_ipd(1)'last_event,  tpd_A_O((511 - 3)- 32*14 ), true),
						5 => (A_ipd(2)'last_event,  tpd_A_O((511 - 3)- 32*13 ), true),
						6 => (A_ipd(3)'last_event,  tpd_A_O((511 - 3)- 32*12 ), true),
						7 => (A_ipd(4)'last_event,  tpd_A_O((511 - 3)- 32*11 ), true), 
						8 => (A_ipd(5)'last_event,  tpd_A_O((511 - 3)- 32*10 ), true),
						9 => (A_ipd(6)'last_event,  tpd_A_O((511 - 3)- 32*9 ), true),
						10 => (A_ipd(7)'last_event,  tpd_A_O((511 - 3)- 32*8 ), true),
						11=> (A_ipd(8)'last_event,  tpd_A_O((511 - 3)- 32*7 ), true),
						12 => (A_ipd(9)'last_event,  tpd_A_O((511 - 3)- 32*6 ), true),
						13 => (A_ipd(10)'last_event,  tpd_A_O((511 - 3)- 32*5 ), true),
						14 => (A_ipd(11)'last_event,  tpd_A_O((511 - 3)- 32*4 ), true),
						15 => (A_ipd(12)'last_event,  tpd_A_O((511 - 3)- 32*3 ), true),
						16=> (A_ipd(13)'last_event,  tpd_A_O((511 - 3)- 32*2), true),
						17=> (A_ipd(14)'last_event,  tpd_A_O((511 - 3)- 32*1 ), true), 
						18=> (A_ipd(15)'last_event,  tpd_A_O((511 - 3)- 32*0 ), true), 
						19=> (B_ipd(0)'last_event,  tpd_B_O((511 - 3)- 32*15 ), true),
						20 => (B_ipd(1)'last_event,  tpd_B_O((511 - 3)- 32*14 ), true),
						21 => (B_ipd(2)'last_event,  tpd_B_O((511 - 3)- 32*13 ), true),
						22 => (B_ipd(3)'last_event,  tpd_B_O((511 - 3)- 32*12 ), true),
						23=> (B_ipd(4)'last_event,  tpd_B_O((511 - 3)- 32*11 ), true), 
						24=> (B_ipd(5)'last_event,  tpd_B_O((511 - 3)- 32*10 ), true),
						25 => (B_ipd(6)'last_event,  tpd_B_O((511 - 3)- 32*9 ), true),
						26 => (B_ipd(7)'last_event,  tpd_B_O((511 - 3)- 32*8 ), true),
						27=> (B_ipd(8)'last_event,  tpd_B_O((511 - 3)- 32*7), true),
						28 => (B_ipd(9)'last_event,  tpd_B_O((511 - 3)- 32*6 ), true),
						29=> (B_ipd(10)'last_event,  tpd_B_O((511 - 3)- 32*5 ), true),
						30 => (B_ipd(11)'last_event,  tpd_B_O((511 - 3)- 32*4 ), true),
						31 => (B_ipd(12)'last_event,  tpd_B_O((511 - 3)- 32*3 ), true),
						32=> (B_ipd(13)'last_event,  tpd_B_O((511 - 3)- 32*2 ), true),
						33=> (B_ipd(14)'last_event,  tpd_B_O((511 - 3)- 32*1 ), true), 
						34=> (B_ipd(15)'last_event,  tpd_B_O((511 - 3)- 32*0 ), true),
						35=> (C_ipd(0)'last_event,  tpd_C_O((511 - 3)- 32*15 ), true),
						36 => (C_ipd(1)'last_event,  tpd_C_O((511 - 3)- 32*14 ), true),
						37 => (C_ipd(2)'last_event,  tpd_C_O((511 - 3)- 32*13 ), true),
						38 => (C_ipd(3)'last_event,  tpd_C_O((511 - 3)- 32*12 ), true),
						39=> (C_ipd(4)'last_event,  tpd_C_O((511 - 3)- 32*11 ), true), 
						40=> (C_ipd(5)'last_event,  tpd_C_O((511 - 3)- 32*10 ), true),
						41 => (C_ipd(6)'last_event,  tpd_C_O((511 - 3)- 32*9 ), true),
						42 => (C_ipd(7)'last_event,  tpd_C_O((511 - 3)- 32*8 ), true),
						43=> (C_ipd(8)'last_event,  tpd_C_O((511 - 3)- 32*7), true),
						44 => (C_ipd(9)'last_event,  tpd_C_O((511 - 3)- 32*6 ), true),
						45=> (C_ipd(10)'last_event,  tpd_C_O((511 - 3)- 32*5 ), true),
						46 => (C_ipd(11)'last_event,  tpd_C_O((511 - 3)- 32*4 ), true),
						47 => (C_ipd(12)'last_event,  tpd_C_O((511 - 3)- 32*3 ), true),
						48=> (C_ipd(13)'last_event,  tpd_C_O((511 - 3)- 32*2 ), true),
						49=> (C_ipd(14)'last_event,  tpd_C_O((511 - 3)- 32*1 ), true), 
						50=> (C_ipd(15)'last_event,  tpd_C_O((511 - 3)- 32*0 ), true),
						51=> (D_ipd(0)'last_event,  tpd_D_O((511 - 3)- 32*15 ), true),
						52 => (D_ipd(1)'last_event,  tpd_D_O((511 - 3)- 32*14 ), true),
						53 => (D_ipd(2)'last_event,  tpd_D_O((511 - 3)- 32*13 ), true),
						54 => (D_ipd(3)'last_event,  tpd_D_O((511 - 3)- 32*12 ), true),
						55=> (D_ipd(4)'last_event,  tpd_D_O((511 - 3)- 32*11 ), true), 
						56=> (D_ipd(5)'last_event,  tpd_D_O((511 - 3)- 32*10 ), true),
						57 => (D_ipd(6)'last_event,  tpd_D_O((511 - 3)- 32*9 ), true),
						58 => (D_ipd(7)'last_event,  tpd_D_O((511 - 3)- 32*8 ), true),
						59=> (D_ipd(8)'last_event,  tpd_D_O((511 - 3)- 32*7 ), true),
						60 => (D_ipd(9)'last_event,  tpd_D_O((511 - 3)- 32*6 ), true),
						61=> (D_ipd(10)'last_event,  tpd_D_O((511 - 3)- 32*5 ), true),
						62 => (D_ipd(11)'last_event,  tpd_D_O((511 - 3)- 32*4 ), true),
						63 => (D_ipd(12)'last_event,  tpd_D_O((511 - 3)- 32*3 ), true),
						64=> (D_ipd(13)'last_event,  tpd_D_O((511 - 3)- 32*2 ), true),
						65=> (D_ipd(14)'last_event,  tpd_D_O((511 - 3)- 32*1 ), true), 
						66=> (D_ipd(15)'last_event,  tpd_D_O((511 - 3)- 32*0 ), true),
						67=> (CI_ipd'last_event, tpd_CI_O(28), true)  ,  
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(28), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(28),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(28),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(28),true)),
      Mode          => VitalTransport,	 
	  IgnoreDefaultDelay => TRUE,	   
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);  
	  
	  
	  
	  	  	  	   VitalPathDelay01 (
      OutSignal     => O(29),
      GlitchData    => O_GlitchData(29),
      OutSignalName => "O(29)",
      OutTemp       => O_zd(29),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(29), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(29), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(29), true),
							3 => (A_ipd(0)'last_event,  tpd_A_O((511 - 2)- 32*15 ), true),
						4 => (A_ipd(1)'last_event,  tpd_A_O((511 - 2)- 32*14 ), true),
						5 => (A_ipd(2)'last_event,  tpd_A_O((511 - 2)- 32*13 ), true),
						6 => (A_ipd(3)'last_event,  tpd_A_O((511 - 2)- 32*12 ), true),
						7 => (A_ipd(4)'last_event,  tpd_A_O((511 - 2)- 32*11 ), true), 
						8 => (A_ipd(5)'last_event,  tpd_A_O((511 - 2)- 32*10 ), true),
						9 => (A_ipd(6)'last_event,  tpd_A_O((511 - 2)- 32*9 ), true),
						10 => (A_ipd(7)'last_event,  tpd_A_O((511 - 2)- 32*8 ), true),
						11=> (A_ipd(8)'last_event,  tpd_A_O((511 - 2)- 32*7 ), true),
						12 => (A_ipd(9)'last_event,  tpd_A_O((511 - 2)- 32*6 ), true),
						13 => (A_ipd(10)'last_event,  tpd_A_O((511 - 2)- 32*5 ), true),
						14 => (A_ipd(11)'last_event,  tpd_A_O((511 - 2)- 32*4 ), true),
						15 => (A_ipd(12)'last_event,  tpd_A_O((511 - 2)- 32*3 ), true),
						16=> (A_ipd(13)'last_event,  tpd_A_O((511 - 2)- 32*2), true),
						17=> (A_ipd(14)'last_event,  tpd_A_O((511 - 2)- 32*1 ), true), 
						18=> (A_ipd(15)'last_event,  tpd_A_O((511 - 2)- 32*0 ), true), 
						19=> (B_ipd(0)'last_event,  tpd_B_O((511 - 2)- 32*15 ), true),
						20 => (B_ipd(1)'last_event,  tpd_B_O((511 - 2)- 32*14 ), true),
						21 => (B_ipd(2)'last_event,  tpd_B_O((511 - 2)- 32*13 ), true),
						22 => (B_ipd(3)'last_event,  tpd_B_O((511 - 2)- 32*12 ), true),
						23=> (B_ipd(4)'last_event,  tpd_B_O((511 - 2)- 32*11 ), true), 
						24=> (B_ipd(5)'last_event,  tpd_B_O((511 - 2)- 32*10 ), true),
						25 => (B_ipd(6)'last_event,  tpd_B_O((511 - 2)- 32*9 ), true),
						26 => (B_ipd(7)'last_event,  tpd_B_O((511 - 2)- 32*8 ), true),
						27=> (B_ipd(8)'last_event,  tpd_B_O((511 - 2)- 32*7), true),
						28 => (B_ipd(9)'last_event,  tpd_B_O((511 - 2)- 32*6 ), true),
						29=> (B_ipd(10)'last_event,  tpd_B_O((511 - 2)- 32*5 ), true),
						30 => (B_ipd(11)'last_event,  tpd_B_O((511 - 2)- 32*4 ), true),
						31 => (B_ipd(12)'last_event,  tpd_B_O((511 - 2)- 32*3 ), true),
						32=> (B_ipd(13)'last_event,  tpd_B_O((511 - 2)- 32*2 ), true),
						33=> (B_ipd(14)'last_event,  tpd_B_O((511 - 2)- 32*1 ), true), 
						34=> (B_ipd(15)'last_event,  tpd_B_O((511 - 2)- 32*0 ), true),
						35=> (C_ipd(0)'last_event,  tpd_C_O((511 - 2)- 32*15 ), true),
						36 => (C_ipd(1)'last_event,  tpd_C_O((511 - 2)- 32*14 ), true),
						37 => (C_ipd(2)'last_event,  tpd_C_O((511 - 2)- 32*13 ), true),
						38 => (C_ipd(3)'last_event,  tpd_C_O((511 - 2)- 32*12 ), true),
						39=> (C_ipd(4)'last_event,  tpd_C_O((511 - 2)- 32*11 ), true), 
						40=> (C_ipd(5)'last_event,  tpd_C_O((511 - 2)- 32*10 ), true),
						41 => (C_ipd(6)'last_event,  tpd_C_O((511 - 2)- 32*9 ), true),
						42 => (C_ipd(7)'last_event,  tpd_C_O((511 - 2)- 32*8 ), true),
						43=> (C_ipd(8)'last_event,  tpd_C_O((511 - 2)- 32*7), true),
						44 => (C_ipd(9)'last_event,  tpd_C_O((511 - 2)- 32*6 ), true),
						45=> (C_ipd(10)'last_event,  tpd_C_O((511 - 2)- 32*5 ), true),
						46 => (C_ipd(11)'last_event,  tpd_C_O((511 - 2)- 32*4 ), true),
						47 => (C_ipd(12)'last_event,  tpd_C_O((511 - 2)- 32*3 ), true),
						48=> (C_ipd(13)'last_event,  tpd_C_O((511 - 2)- 32*2 ), true),
						49=> (C_ipd(14)'last_event,  tpd_C_O((511 - 2)- 32*1 ), true), 
						50=> (C_ipd(15)'last_event,  tpd_C_O((511 - 2)- 32*0 ), true),
						51=> (D_ipd(0)'last_event,  tpd_D_O((511 - 2)- 32*15 ), true),
						52 => (D_ipd(1)'last_event,  tpd_D_O((511 - 2)- 32*14 ), true),
						53 => (D_ipd(2)'last_event,  tpd_D_O((511 - 2)- 32*13 ), true),
						54 => (D_ipd(3)'last_event,  tpd_D_O((511 - 2)- 32*12 ), true),
						55=> (D_ipd(4)'last_event,  tpd_D_O((511 - 2)- 32*11 ), true), 
						56=> (D_ipd(5)'last_event,  tpd_D_O((511 - 2)- 32*10 ), true),
						57 => (D_ipd(6)'last_event,  tpd_D_O((511 - 2)- 32*9 ), true),
						58 => (D_ipd(7)'last_event,  tpd_D_O((511 - 2)- 32*8 ), true),
						59=> (D_ipd(8)'last_event,  tpd_D_O((511 - 2)- 32*7 ), true),
						60 => (D_ipd(9)'last_event,  tpd_D_O((511 - 2)- 32*6 ), true),
						61=> (D_ipd(10)'last_event,  tpd_D_O((511 - 2)- 32*5 ), true),
						62 => (D_ipd(11)'last_event,  tpd_D_O((511 - 2)- 32*4 ), true),
						63 => (D_ipd(12)'last_event,  tpd_D_O((511 - 2)- 32*3 ), true),
						64=> (D_ipd(13)'last_event,  tpd_D_O((511 - 2)- 32*2 ), true),
						65=> (D_ipd(14)'last_event,  tpd_D_O((511 - 2)- 32*1 ), true), 
						66=> (D_ipd(15)'last_event,  tpd_D_O((511 - 2)- 32*0 ), true),
						67=> (CI_ipd'last_event, tpd_CI_O(29), true)  ,  
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(29), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(29),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(29),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(29),true)),
      Mode          => VitalTransport,		
	  IgnoreDefaultDelay => TRUE,	 
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);  	
	  
	  
	  
	  	  	  	   VitalPathDelay01 (
      OutSignal     => O(30),
      GlitchData    => O_GlitchData(30),
      OutSignalName => "O(30)",
      OutTemp       => O_zd(30),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(30), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(30), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(30), true),
							3 => (A_ipd(0)'last_event,  tpd_A_O((511 - 1)- 32*15 ), true),
						4 => (A_ipd(1)'last_event,  tpd_A_O((511 - 1)- 32*14 ), true),
						5 => (A_ipd(2)'last_event,  tpd_A_O((511 - 1)- 32*13 ), true),
						6 => (A_ipd(3)'last_event,  tpd_A_O((511 - 1)- 32*12 ), true),
						7 => (A_ipd(4)'last_event,  tpd_A_O((511 - 1)- 32*11 ), true), 
						8 => (A_ipd(5)'last_event,  tpd_A_O((511 - 1)- 32*10 ), true),
						9 => (A_ipd(6)'last_event,  tpd_A_O((511 - 1)- 32*9 ), true),
						10 => (A_ipd(7)'last_event,  tpd_A_O((511 - 1)- 32*8 ), true),
						11=> (A_ipd(8)'last_event,  tpd_A_O((511 - 1)- 32*7 ), true),
						12 => (A_ipd(9)'last_event,  tpd_A_O((511 - 1)- 32*6 ), true),
						13 => (A_ipd(10)'last_event,  tpd_A_O((511 - 1)- 32*5 ), true),
						14 => (A_ipd(11)'last_event,  tpd_A_O((511 - 1)- 32*4 ), true),
						15 => (A_ipd(12)'last_event,  tpd_A_O((511 - 1)- 32*3 ), true),
						16=> (A_ipd(13)'last_event,  tpd_A_O((511 - 1)- 32*2), true),
						17=> (A_ipd(14)'last_event,  tpd_A_O((511 - 1)- 32*1 ), true), 
						18=> (A_ipd(15)'last_event,  tpd_A_O((511 - 1)- 32*0 ), true), 
						19=> (B_ipd(0)'last_event,  tpd_B_O((511 - 1)- 32*15 ), true),
						20 => (B_ipd(1)'last_event,  tpd_B_O((511 - 1)- 32*14 ), true),
						21 => (B_ipd(2)'last_event,  tpd_B_O((511 - 1)- 32*13 ), true),
						22 => (B_ipd(3)'last_event,  tpd_B_O((511 - 1)- 32*12 ), true),
						23=> (B_ipd(4)'last_event,  tpd_B_O((511 - 1)- 32*11 ), true), 
						24=> (B_ipd(5)'last_event,  tpd_B_O((511 - 1)- 32*10 ), true),
						25 => (B_ipd(6)'last_event,  tpd_B_O((511 - 1)- 32*9 ), true),
						26 => (B_ipd(7)'last_event,  tpd_B_O((511 - 1)- 32*8 ), true),
						27=> (B_ipd(8)'last_event,  tpd_B_O((511 - 1)- 32*7), true),
						28 => (B_ipd(9)'last_event,  tpd_B_O((511 - 1)- 32*6 ), true),
						29=> (B_ipd(10)'last_event,  tpd_B_O((511 - 1)- 32*5 ), true),
						30 => (B_ipd(11)'last_event,  tpd_B_O((511 - 1)- 32*4 ), true),
						31 => (B_ipd(12)'last_event,  tpd_B_O((511 - 1)- 32*3 ), true),
						32=> (B_ipd(13)'last_event,  tpd_B_O((511 - 1)- 32*2 ), true),
						33=> (B_ipd(14)'last_event,  tpd_B_O((511 - 1)- 32*1 ), true), 
						34=> (B_ipd(15)'last_event,  tpd_B_O((511 - 1)- 32*0 ), true),
						35=> (C_ipd(0)'last_event,  tpd_C_O((511 - 1)- 32*15 ), true),
						36 => (C_ipd(1)'last_event,  tpd_C_O((511 - 1)- 32*14 ), true),
						37 => (C_ipd(2)'last_event,  tpd_C_O((511 - 1)- 32*13 ), true),
						38 => (C_ipd(3)'last_event,  tpd_C_O((511 - 1)- 32*12 ), true),
						39=> (C_ipd(4)'last_event,  tpd_C_O((511 - 1)- 32*11 ), true), 
						40=> (C_ipd(5)'last_event,  tpd_C_O((511 - 1)- 32*10 ), true),
						41 => (C_ipd(6)'last_event,  tpd_C_O((511 - 1)- 32*9 ), true),
						42 => (C_ipd(7)'last_event,  tpd_C_O((511 - 1)- 32*8 ), true),
						43=> (C_ipd(8)'last_event,  tpd_C_O((511 - 1)- 32*7), true),
						44 => (C_ipd(9)'last_event,  tpd_C_O((511 - 1)- 32*6 ), true),
						45=> (C_ipd(10)'last_event,  tpd_C_O((511 - 1)- 32*5 ), true),
						46 => (C_ipd(11)'last_event,  tpd_C_O((511 - 1)- 32*4 ), true),
						47 => (C_ipd(12)'last_event,  tpd_C_O((511 - 1)- 32*3 ), true),
						48=> (C_ipd(13)'last_event,  tpd_C_O((511 - 1)- 32*2 ), true),
						49=> (C_ipd(14)'last_event,  tpd_C_O((511 - 1)- 32*1 ), true), 
						50=> (C_ipd(15)'last_event,  tpd_C_O((511 - 1)- 32*0 ), true),
						51=> (D_ipd(0)'last_event,  tpd_D_O((511 - 1)- 32*15 ), true),
						52 => (D_ipd(1)'last_event,  tpd_D_O((511 - 1)- 32*14 ), true),
						53 => (D_ipd(2)'last_event,  tpd_D_O((511 - 1)- 32*13 ), true),
						54 => (D_ipd(3)'last_event,  tpd_D_O((511 - 1)- 32*12 ), true),
						55=> (D_ipd(4)'last_event,  tpd_D_O((511 - 1)- 32*11 ), true), 
						56=> (D_ipd(5)'last_event,  tpd_D_O((511 - 1)- 32*10 ), true),
						57 => (D_ipd(6)'last_event,  tpd_D_O((511 - 1)- 32*9 ), true),
						58 => (D_ipd(7)'last_event,  tpd_D_O((511 - 1)- 32*8 ), true),
						59=> (D_ipd(8)'last_event,  tpd_D_O((511 - 1)- 32*7 ), true),
						60 => (D_ipd(9)'last_event,  tpd_D_O((511 - 1)- 32*6 ), true),
						61=> (D_ipd(10)'last_event,  tpd_D_O((511 - 1)- 32*5 ), true),
						62 => (D_ipd(11)'last_event,  tpd_D_O((511 - 1)- 32*4 ), true),
						63 => (D_ipd(12)'last_event,  tpd_D_O((511 - 1)- 32*3 ), true),
						64=> (D_ipd(13)'last_event,  tpd_D_O((511 - 1)- 32*2 ), true),
						65=> (D_ipd(14)'last_event,  tpd_D_O((511 - 1)- 32*1 ), true), 
						66=> (D_ipd(15)'last_event,  tpd_D_O((511 - 1)- 32*0 ), true),
						67=> (CI_ipd'last_event, tpd_CI_O(30), true) ,  
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(30), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(30),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(30),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(30),true)),
      Mode          => VitalTransport,		  
	  IgnoreDefaultDelay => TRUE,		  
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);  	  
	  
	  
	  	  	  	   VitalPathDelay01 (
      OutSignal     => O(31),
      GlitchData    => O_GlitchData(31),
      OutSignalName => "O(31)",
      OutTemp       => O_zd(31),
      Paths         => (0 => (CLK_ipd'last_event, tpd_CLK_O_posedge(31), true),
	  					1 => (ORSTBOT_ipd'last_event, tpd_ORSTBOT_O(31), true),
	  					2 => (ORSTTOP_ipd'last_event, tpd_ORSTTOP_O(31), true),
							3 => (A_ipd(0)'last_event,  tpd_A_O((511 - 0)- 32*15 ), true),
						4 => (A_ipd(1)'last_event,  tpd_A_O((511 - 0)- 32*14 ), true),
						5 => (A_ipd(2)'last_event,  tpd_A_O((511 - 0)- 32*13 ), true),
						6 => (A_ipd(3)'last_event,  tpd_A_O((511 - 0)- 32*12 ), true),
						7 => (A_ipd(4)'last_event,  tpd_A_O((511 - 0)- 32*11 ), true), 
						8 => (A_ipd(5)'last_event,  tpd_A_O((511 - 0)- 32*10 ), true),
						9 => (A_ipd(6)'last_event,  tpd_A_O((511 - 0)- 32*9 ), true),
						10 => (A_ipd(7)'last_event,  tpd_A_O((511 - 0)- 32*8 ), true),
						11=> (A_ipd(8)'last_event,  tpd_A_O((511 - 0)- 32*7 ), true),
						12 => (A_ipd(9)'last_event,  tpd_A_O((511 - 0)- 32*6 ), true),
						13 => (A_ipd(10)'last_event,  tpd_A_O((511 - 0)- 32*5 ), true),
						14 => (A_ipd(11)'last_event,  tpd_A_O((511 - 0)- 32*4 ), true),
						15 => (A_ipd(12)'last_event,  tpd_A_O((511 - 0)- 32*3 ), true),
						16=> (A_ipd(13)'last_event,  tpd_A_O((511 - 0)- 32*2), true),
						17=> (A_ipd(14)'last_event,  tpd_A_O((511 - 0)- 32*1 ), true), 
						18=> (A_ipd(15)'last_event,  tpd_A_O((511 - 0)- 32*0 ), true), 
						19=> (B_ipd(0)'last_event,  tpd_B_O((511 - 0)- 32*15 ), true),
						20 => (B_ipd(1)'last_event,  tpd_B_O((511 - 0)- 32*14 ), true),
						21 => (B_ipd(2)'last_event,  tpd_B_O((511 - 0)- 32*13 ), true),
						22 => (B_ipd(3)'last_event,  tpd_B_O((511 - 0)- 32*12 ), true),
						23=> (B_ipd(4)'last_event,  tpd_B_O((511 - 0)- 32*11 ), true), 
						24=> (B_ipd(5)'last_event,  tpd_B_O((511 - 0)- 32*10 ), true),
						25 => (B_ipd(6)'last_event,  tpd_B_O((511 - 0)- 32*9 ), true),
						26 => (B_ipd(7)'last_event,  tpd_B_O((511 - 0)- 32*8 ), true),
						27=> (B_ipd(8)'last_event,  tpd_B_O((511 - 0)- 32*7), true),
						28 => (B_ipd(9)'last_event,  tpd_B_O((511 - 0)- 32*6 ), true),
						29=> (B_ipd(10)'last_event,  tpd_B_O((511 - 0)- 32*5 ), true),
						30 => (B_ipd(11)'last_event,  tpd_B_O((511 - 0)- 32*4 ), true),
						31 => (B_ipd(12)'last_event,  tpd_B_O((511 - 0)- 32*3 ), true),
						32=> (B_ipd(13)'last_event,  tpd_B_O((511 - 0)- 32*2 ), true),
						33=> (B_ipd(14)'last_event,  tpd_B_O((511 - 0)- 32*1 ), true), 
						34=> (B_ipd(15)'last_event,  tpd_B_O((511 - 0)- 32*0 ), true),
						35=> (C_ipd(0)'last_event,  tpd_C_O((511 - 0)- 32*15 ), true),
						36 => (C_ipd(1)'last_event,  tpd_C_O((511 - 0)- 32*14 ), true),
						37 => (C_ipd(2)'last_event,  tpd_C_O((511 - 0)- 32*13 ), true),
						38 => (C_ipd(3)'last_event,  tpd_C_O((511 - 0)- 32*12 ), true),
						39=> (C_ipd(4)'last_event,  tpd_C_O((511 - 0)- 32*11 ), true), 
						40=> (C_ipd(5)'last_event,  tpd_C_O((511 - 0)- 32*10 ), true),
						41 => (C_ipd(6)'last_event,  tpd_C_O((511 - 0)- 32*9 ), true),
						42 => (C_ipd(7)'last_event,  tpd_C_O((511 - 0)- 32*8 ), true),
						43=> (C_ipd(8)'last_event,  tpd_C_O((511 - 0)- 32*7), true),
						44 => (C_ipd(9)'last_event,  tpd_C_O((511 - 0)- 32*6 ), true),
						45=> (C_ipd(10)'last_event,  tpd_C_O((511 - 0)- 32*5 ), true),
						46 => (C_ipd(11)'last_event,  tpd_C_O((511 - 0)- 32*4 ), true),
						47 => (C_ipd(12)'last_event,  tpd_C_O((511 - 0)- 32*3 ), true),
						48=> (C_ipd(13)'last_event,  tpd_C_O((511 - 0)- 32*2 ), true),
						49=> (C_ipd(14)'last_event,  tpd_C_O((511 - 0)- 32*1 ), true), 
						50=> (C_ipd(15)'last_event,  tpd_C_O((511 - 0)- 32*0 ), true),
						51=> (D_ipd(0)'last_event,  tpd_D_O((511 - 0)- 32*15 ), true),
						52 => (D_ipd(1)'last_event,  tpd_D_O((511 - 0)- 32*14 ), true),
						53 => (D_ipd(2)'last_event,  tpd_D_O((511 - 0)- 32*13 ), true),
						54 => (D_ipd(3)'last_event,  tpd_D_O((511 - 0)- 32*12 ), true),
						55=> (D_ipd(4)'last_event,  tpd_D_O((511 - 0)- 32*11 ), true), 
						56=> (D_ipd(5)'last_event,  tpd_D_O((511 - 0)- 32*10 ), true),
						57 => (D_ipd(6)'last_event,  tpd_D_O((511 - 0)- 32*9 ), true),
						58 => (D_ipd(7)'last_event,  tpd_D_O((511 - 0)- 32*8 ), true),
						59=> (D_ipd(8)'last_event,  tpd_D_O((511 - 0)- 32*7 ), true),
						60 => (D_ipd(9)'last_event,  tpd_D_O((511 - 0)- 32*6 ), true),
						61=> (D_ipd(10)'last_event,  tpd_D_O((511 - 0)- 32*5 ), true),
						62 => (D_ipd(11)'last_event,  tpd_D_O((511 - 0)- 32*4 ), true),
						63 => (D_ipd(12)'last_event,  tpd_D_O((511 - 0)- 32*3 ), true),
						64=> (D_ipd(13)'last_event,  tpd_D_O((511 - 0)- 32*2 ), true),
						65=> (D_ipd(14)'last_event,  tpd_D_O((511 - 0)- 32*1 ), true), 
						66=> (D_ipd(15)'last_event,  tpd_D_O((511 - 0)- 32*0 ), true),
						67=> (CI_ipd'last_event, tpd_CI_O(31), true)  ,  
						68=> (ADDSUBTOP_ipd'last_event,  tpd_ADDSUBTOP_O(31), true),
						69=> (ADDSUBBOT_ipd'last_event,tpd_ADDSUBBOT_O(31),true),
					   	70=>  (OLOADTOP_ipd'last_event,tpd_OLOADTOP_O(31),true),	 
						71=>  (OLOADBOT_ipd'last_event,tpd_OLOADBOT_O(31),true)),
      Mode          => VitalTransport,					
	  IgnoreDefaultDelay => TRUE,						  
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);  
	  
	  
	  
	  	  	  	   VitalPathDelay01 (
      OutSignal     => CO,
      GlitchData    => CO_GlitchData,
      OutSignalName => "CO",
      OutTemp       => CO_zd,
      Paths         => (0 => (A_ipd(0)'last_event,  tpd_A_CO(0), true),
						1 => (A_ipd(1)'last_event,  tpd_A_CO(1), true),
						2 => (A_ipd(2)'last_event,  tpd_A_CO(2), true),
						3 => (A_ipd(3)'last_event,  tpd_A_CO(3), true),
						4 => (A_ipd(4)'last_event,  tpd_A_CO(4), true), 
						5 => (A_ipd(5)'last_event,  tpd_A_CO(5), true),
						6 => (A_ipd(6)'last_event,  tpd_A_CO(6), true),
						7 => (A_ipd(7)'last_event,  tpd_A_CO(7), true),
						8=> (A_ipd(8)'last_event,  tpd_A_CO(8 ), true),
						9 => (A_ipd(9)'last_event,  tpd_A_CO(9), true),
						10 => (A_ipd(10)'last_event,  tpd_A_CO(10 ), true),
						11 => (A_ipd(11)'last_event,  tpd_A_CO(11), true),
						12 => (A_ipd(12)'last_event,  tpd_A_CO(12 ), true),
						13=> (A_ipd(13)'last_event,  tpd_A_CO(13), true),
						14=> (A_ipd(14)'last_event,  tpd_A_CO(14), true), 
						15=> (A_ipd(15)'last_event,  tpd_A_CO(15 ), true)
						),
      Mode          => VitalTransport,					
	  IgnoreDefaultDelay => TRUE,						  
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning); 		
	  
	    	  	  	   VitalPathDelay01 (
      OutSignal     => CO,
      GlitchData    => CO_GlitchData,
      OutSignalName => "CO",
      OutTemp       => CO_zd,
      Paths         => (0 => (B_ipd(0)'last_event,  tpd_B_CO(0), true),
						1 => (B_ipd(1)'last_event,  tpd_B_CO(1), true),
						2 => (B_ipd(2)'last_event,  tpd_B_CO(2), true),
						3 => (B_ipd(3)'last_event,  tpd_B_CO(3), true),
						4 => (B_ipd(4)'last_event,  tpd_B_CO(4), true), 
						5 => (B_ipd(5)'last_event,  tpd_B_CO(5), true),
						6 => (B_ipd(6)'last_event,  tpd_B_CO(6), true),
						7 => (B_ipd(7)'last_event,  tpd_B_CO(7), true),
						8=> (B_ipd(8)'last_event,  tpd_B_CO(8 ), true),
						9 => (B_ipd(9)'last_event,  tpd_B_CO(9), true),
						10 => (B_ipd(10)'last_event,  tpd_B_CO(10 ), true),
						11 => (B_ipd(11)'last_event,  tpd_B_CO(11), true),
						12 => (B_ipd(12)'last_event,  tpd_B_CO(12 ), true),
						13=> (B_ipd(13)'last_event,  tpd_B_CO(13), true),
						14=> (B_ipd(14)'last_event,  tpd_B_CO(14), true), 
						15=> (B_ipd(15)'last_event,  tpd_B_CO(15 ), true)
						),
      Mode          => VitalTransport,					
	  IgnoreDefaultDelay => TRUE,						  
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning); 
	  
	    	  	  	   VitalPathDelay01 (
      OutSignal     => CO,
      GlitchData    => CO_GlitchData,
      OutSignalName => "CO",
      OutTemp       => CO_zd,
      Paths         => (0 => (C_ipd(0)'last_event,  tpd_C_CO(0), true),
						1 => (C_ipd(1)'last_event,  tpd_C_CO(1), true),
						2 => (C_ipd(2)'last_event,  tpd_C_CO(2), true),
						3 => (C_ipd(3)'last_event,  tpd_C_CO(3), true),
						4 => (C_ipd(4)'last_event,  tpd_C_CO(4), true), 
						5 => (C_ipd(5)'last_event,  tpd_C_CO(5), true),
						6 => (C_ipd(6)'last_event,  tpd_C_CO(6), true),
						7 => (C_ipd(7)'last_event,  tpd_C_CO(7), true),
						8=> (C_ipd(8)'last_event,  tpd_C_CO(8 ), true),
						9 => (C_ipd(9)'last_event,  tpd_C_CO(9), true),
						10 => (C_ipd(10)'last_event,  tpd_C_CO(10 ), true),
						11 => (C_ipd(11)'last_event,  tpd_C_CO(11), true),
						12 => (C_ipd(12)'last_event,  tpd_C_CO(12 ), true),
						13=> (C_ipd(13)'last_event,  tpd_C_CO(13), true),
						14=> (C_ipd(14)'last_event,  tpd_C_CO(14), true), 
						15=> (C_ipd(15)'last_event,  tpd_C_CO(15 ), true)
						),
      Mode          => VitalTransport,					
	  IgnoreDefaultDelay => TRUE,						  
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning); 
	  
	  
	    	  	  	   VitalPathDelay01 (
      OutSignal     => CO,
      GlitchData    => CO_GlitchData,
      OutSignalName => "CO",
      OutTemp       => CO_zd,
      Paths         => (0 => (D_ipd(0)'last_event,  tpd_D_CO(0), true),
						1 => (D_ipd(1)'last_event,  tpd_D_CO(1), true),
						2 => (D_ipd(2)'last_event,  tpd_D_CO(2), true),
						3 => (D_ipd(3)'last_event,  tpd_D_CO(3), true),
						4 => (D_ipd(4)'last_event,  tpd_D_CO(4), true), 
						5 => (D_ipd(5)'last_event,  tpd_D_CO(5), true),
						6 => (D_ipd(6)'last_event,  tpd_D_CO(6), true),
						7 => (D_ipd(7)'last_event,  tpd_D_CO(7), true),
						8=> (D_ipd(8)'last_event,  tpd_D_CO(8 ), true),
						9 => (D_ipd(9)'last_event,  tpd_D_CO(9), true),
						10 => (D_ipd(10)'last_event,  tpd_D_CO(10 ), true),
						11 => (D_ipd(11)'last_event,  tpd_D_CO(11), true),
						12 => (D_ipd(12)'last_event,  tpd_D_CO(12 ), true),
						13=> (D_ipd(13)'last_event,  tpd_D_CO(13), true),
						14=> (D_ipd(14)'last_event,  tpd_D_CO(14), true), 
						15=> (D_ipd(15)'last_event,  tpd_D_CO(15 ), true)
						),
      Mode          => VitalTransport,					
	  IgnoreDefaultDelay => TRUE,						  
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning); 
	  
	  
	  
	    	  	  	   VitalPathDelay01 (
      OutSignal     => CO,
      GlitchData    => CO_GlitchData,
      OutSignalName => "CO",
      OutTemp       => CO_zd,
      Paths         => (0 => (CI_ipd'last_event,  tpd_CI_CO, true)
						),
      Mode          => VitalTransport,					
	  IgnoreDefaultDelay => TRUE,						  
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);


  	  	  	   VitalPathDelay01 (
      OutSignal     => CO,
      GlitchData    => CO_GlitchData,
      OutSignalName => "CO",
      OutTemp       => CO_zd,
      Paths         => (0 => (ACCUMCI_ipd'last_event,  tpd_ACCUMCI_CO, true)
						),
      Mode          => VitalTransport,					
	  IgnoreDefaultDelay => TRUE,						  
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning); 	  
	  
	  
	    	  	  	   VitalPathDelay01 (
      OutSignal     => CO,
      GlitchData    => CO_GlitchData,
      OutSignalName => "CO",
      OutTemp       => CO_zd,
      Paths         => (0 => (CLK_ipd'last_event,  tpd_CLK_CO_posedge, true)
						),
      Mode          => VitalTransport,					
	  IgnoreDefaultDelay => TRUE,						  
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning); 
	  
	  
	    	  	  	   VitalPathDelay01 (
      OutSignal     => CO,
      GlitchData    => CO_GlitchData,
      OutSignalName => "CO",
      OutTemp       => CO_zd,
      Paths         => (0 => (ADDSUBBOT_ipd'last_event,  tpd_ADDSUBBOT_CO, true)
						),
      Mode          => VitalTransport,					
	  IgnoreDefaultDelay => TRUE,						  
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning); 
	  
	  
	    	  	  	   VitalPathDelay01 (
      OutSignal     => CO,
      GlitchData    => CO_GlitchData,
      OutSignalName => "CO",
      OutTemp       => CO_zd,
      Paths         => (0 => (OLOADBOT_ipd'last_event,  tpd_OLOADBOT_CO, true)
						),
      Mode          => VitalTransport,					
	  IgnoreDefaultDelay => TRUE,						  
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning); 
	  
	    	  	  	   VitalPathDelay01 (
      OutSignal     => CO,
      GlitchData    => CO_GlitchData,
      OutSignalName => "CO",
      OutTemp       => CO_zd,
      Paths         => (0 => (OLOADTOP_ipd'last_event,  tpd_OLOADTOP_CO, true)),
      Mode          => VitalTransport,					
	  IgnoreDefaultDelay => TRUE,						  
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning); 
	  
	    VitalPathDelay01 (
      OutSignal     => ACCUMCO,
      GlitchData    => ACCUMCO_GlitchData,
      OutSignalName => "ACCUMCO",
      OutTemp       => ACCUMCO_zd,
      Paths         => (0 => (A_ipd(0)'last_event,  tpd_A_ACCUMCO(0), true),
						1 => (A_ipd(1)'last_event,  tpd_A_ACCUMCO(1), true),
						2 => (A_ipd(2)'last_event,  tpd_A_ACCUMCO(2), true),
						3 => (A_ipd(3)'last_event,  tpd_A_ACCUMCO(3), true),
						4 => (A_ipd(4)'last_event,  tpd_A_ACCUMCO(4), true), 
						5 => (A_ipd(5)'last_event,  tpd_A_ACCUMCO(5), true),
						6 => (A_ipd(6)'last_event,  tpd_A_ACCUMCO(6), true),
						7 => (A_ipd(7)'last_event,  tpd_A_ACCUMCO(7), true),
						8=> (A_ipd(8)'last_event,  tpd_A_ACCUMCO(8 ), true),
						9 => (A_ipd(9)'last_event,  tpd_A_ACCUMCO(9), true),
						10 => (A_ipd(10)'last_event,  tpd_A_ACCUMCO(10 ), true),
						11 => (A_ipd(11)'last_event,  tpd_A_ACCUMCO(11), true),
						12 => (A_ipd(12)'last_event,  tpd_A_ACCUMCO(12 ), true),
						13=> (A_ipd(13)'last_event,  tpd_A_ACCUMCO(13), true),
						14=> (A_ipd(14)'last_event,  tpd_A_ACCUMCO(14), true), 
						15=> (A_ipd(15)'last_event,  tpd_A_ACCUMCO(15 ), true)
						),
      Mode          => VitalTransport,					
	  IgnoreDefaultDelay => TRUE,						  
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning); 
	  
	  
	  	    	  	  	   VitalPathDelay01 (
      OutSignal     => ACCUMCO,
      GlitchData    => ACCUMCO_GlitchData,
      OutSignalName => "ACCUMCO",
      OutTemp       => ACCUMCO_zd,
      Paths         => (0 => (B_ipd(0)'last_event,  tpd_B_ACCUMCO(0), true),
						1 => (B_ipd(1)'last_event,  tpd_B_ACCUMCO(1), true),
						2 => (B_ipd(2)'last_event,  tpd_B_ACCUMCO(2), true),
						3 => (B_ipd(3)'last_event,  tpd_B_ACCUMCO(3), true),
						4 => (B_ipd(4)'last_event,  tpd_B_ACCUMCO(4), true), 
						5 => (B_ipd(5)'last_event,  tpd_B_ACCUMCO(5), true),
						6 => (B_ipd(6)'last_event,  tpd_B_ACCUMCO(6), true),
						7 => (B_ipd(7)'last_event,  tpd_B_ACCUMCO(7), true),
						8=> (B_ipd(8)'last_event,  tpd_B_ACCUMCO(8 ), true),
						9 => (B_ipd(9)'last_event,  tpd_B_ACCUMCO(9), true),
						10 => (B_ipd(10)'last_event,  tpd_B_ACCUMCO(10 ), true),
						11 => (B_ipd(11)'last_event,  tpd_B_ACCUMCO(11), true),
						12 => (B_ipd(12)'last_event,  tpd_B_ACCUMCO(12 ), true),
						13=> (B_ipd(13)'last_event,  tpd_B_ACCUMCO(13), true),
						14=> (B_ipd(14)'last_event,  tpd_B_ACCUMCO(14), true), 
						15=> (B_ipd(15)'last_event,  tpd_B_ACCUMCO(15 ), true)
						),
      Mode          => VitalTransport,					
	  IgnoreDefaultDelay => TRUE,						  
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning); 
	  
	    	  	  	   VitalPathDelay01 (
      OutSignal     => ACCUMCO,
      GlitchData    => ACCUMCO_GlitchData,
      OutSignalName => "ACCUMCO",
      OutTemp       => ACCUMCO_zd,
      Paths         => (0 => (C_ipd(0)'last_event,  tpd_C_ACCUMCO(0), true),
						1 => (C_ipd(1)'last_event,  tpd_C_ACCUMCO(1), true),
						2 => (C_ipd(2)'last_event,  tpd_C_ACCUMCO(2), true),
						3 => (C_ipd(3)'last_event,  tpd_C_ACCUMCO(3), true),
						4 => (C_ipd(4)'last_event,  tpd_C_ACCUMCO(4), true), 
						5 => (C_ipd(5)'last_event,  tpd_C_ACCUMCO(5), true),
						6 => (C_ipd(6)'last_event,  tpd_C_ACCUMCO(6), true),
						7 => (C_ipd(7)'last_event,  tpd_C_ACCUMCO(7), true),
						8=> (C_ipd(8)'last_event,  tpd_C_ACCUMCO(8 ), true),
						9 => (C_ipd(9)'last_event,  tpd_C_ACCUMCO(9), true),
						10 => (C_ipd(10)'last_event,  tpd_C_ACCUMCO(10 ), true),
						11 => (C_ipd(11)'last_event,  tpd_C_ACCUMCO(11), true),
						12 => (C_ipd(12)'last_event,  tpd_C_ACCUMCO(12 ), true),
						13=> (C_ipd(13)'last_event,  tpd_C_ACCUMCO(13), true),
						14=> (C_ipd(14)'last_event,  tpd_C_ACCUMCO(14), true), 
						15=> (C_ipd(15)'last_event,  tpd_C_ACCUMCO(15 ), true)
						),
      Mode          => VitalTransport,					
	  IgnoreDefaultDelay => TRUE,						  
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning); 
	  
	  
	    	  	  	   VitalPathDelay01 (
      OutSignal     => ACCUMCO,
      GlitchData    => ACCUMCO_GlitchData,
      OutSignalName => "ACCUMCO",
      OutTemp       => ACCUMCO_zd,
      Paths         => (0 => (D_ipd(0)'last_event,  tpd_D_ACCUMCO(0), true),
						1 => (D_ipd(1)'last_event,  tpd_D_ACCUMCO(1), true),
						2 => (D_ipd(2)'last_event,  tpd_D_ACCUMCO(2), true),
						3 => (D_ipd(3)'last_event,  tpd_D_ACCUMCO(3), true),
						4 => (D_ipd(4)'last_event,  tpd_D_ACCUMCO(4), true), 
						5 => (D_ipd(5)'last_event,  tpd_D_ACCUMCO(5), true),
						6 => (D_ipd(6)'last_event,  tpd_D_ACCUMCO(6), true),
						7 => (D_ipd(7)'last_event,  tpd_D_ACCUMCO(7), true),
						8=> (D_ipd(8)'last_event,  tpd_D_ACCUMCO(8 ), true),
						9 => (D_ipd(9)'last_event,  tpd_D_ACCUMCO(9), true),
						10 => (D_ipd(10)'last_event,  tpd_D_ACCUMCO(10 ), true),
						11 => (D_ipd(11)'last_event,  tpd_D_ACCUMCO(11), true),
						12 => (D_ipd(12)'last_event,  tpd_D_ACCUMCO(12 ), true),
						13=> (D_ipd(13)'last_event,  tpd_D_ACCUMCO(13), true),
						14=> (D_ipd(14)'last_event,  tpd_D_ACCUMCO(14), true), 
						15=> (D_ipd(15)'last_event,  tpd_D_ACCUMCO(15 ), true)
						),
      Mode          => VitalTransport,					
	  IgnoreDefaultDelay => TRUE,						  
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning); 
	  
	  
	  
	    	  	  	   VitalPathDelay01 (
      OutSignal     => ACCUMCO,
      GlitchData    => ACCUMCO_GlitchData,
      OutSignalName => "ACCUMCO",
      OutTemp       => ACCUMCO_zd,
      Paths         => (0 => (CI_ipd'last_event,  tpd_CI_ACCUMCO, true)
						),
      Mode          => VitalTransport,					
	  IgnoreDefaultDelay => TRUE,						  
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);


  	  	  	   VitalPathDelay01 (
      OutSignal     => ACCUMCO,
      GlitchData    => ACCUMCO_GlitchData,
      OutSignalName => "ACCUMCO",
      OutTemp       => ACCUMCO_zd,
      Paths         => (0 => (ACCUMCI_ipd'last_event,  tpd_ACCUMCI_ACCUMCO, true)
						),
      Mode          => VitalTransport,					
	  IgnoreDefaultDelay => TRUE,						  
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning); 	  
	  
	  
	    	  	  	   VitalPathDelay01 (
      OutSignal     => ACCUMCO,
      GlitchData    => ACCUMCO_GlitchData,
      OutSignalName => "ACCUMCO",
      OutTemp       => ACCUMCO_zd,
      Paths         => (0 => (CLK_ipd'last_event,  tpd_CLK_ACCUMCO_posedge, true)
						),
      Mode          => VitalTransport,					
	  IgnoreDefaultDelay => TRUE,						  
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning); 
	  
	  
	    	  	  	   VitalPathDelay01 (
      OutSignal     => ACCUMCO,
      GlitchData    => ACCUMCO_GlitchData,
      OutSignalName => "ACCUMCO",
      OutTemp       => ACCUMCO_zd,
      Paths         => (0 => (ADDSUBBOT_ipd'last_event,  tpd_ADDSUBBOT_ACCUMCO, true)
						),
      Mode          => VitalTransport,					
	  IgnoreDefaultDelay => TRUE,						  
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning); 
	  
	  
	    	  	  	   VitalPathDelay01 (
      OutSignal     => ACCUMCO,
      GlitchData    => ACCUMCO_GlitchData,
      OutSignalName => "ACCUMCO",
      OutTemp       => ACCUMCO_zd,
      Paths         => (0 => (OLOADBOT_ipd'last_event,  tpd_OLOADBOT_ACCUMCO, true)
						),
      Mode          => VitalTransport,					
	  IgnoreDefaultDelay => TRUE,						  
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning); 
	  
	    	  	  	   VitalPathDelay01 (
      OutSignal     => ACCUMCO,
      GlitchData    => ACCUMCO_GlitchData,
      OutSignalName => "ACCUMCO",
      OutTemp       => ACCUMCO_zd,
      Paths         => (0 => (OLOADTOP_ipd'last_event,  tpd_OLOADTOP_ACCUMCO, true)
						),
      Mode          => VitalTransport,					
	  IgnoreDefaultDelay => TRUE,						  
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning); 
	  
	   VitalPathDelay01 (
      OutSignal     => SIGNEXTOUT,
      GlitchData    => SIGNEXTOUT_GlitchData,
      OutSignalName => "SIGNEXTOUT",
      OutTemp       => SIGNEXTOUT_zd,
      Paths         => (0 => (A_ipd(0)'last_event,  tpd_A_SIGNEXTOUT(0), true),
						1 => (A_ipd(1)'last_event,  tpd_A_SIGNEXTOUT(1), true),
						2 => (A_ipd(2)'last_event,  tpd_A_SIGNEXTOUT(2), true),
						3 => (A_ipd(3)'last_event,  tpd_A_SIGNEXTOUT(3), true),
						4 => (A_ipd(4)'last_event,  tpd_A_SIGNEXTOUT(4), true), 
						5 => (A_ipd(5)'last_event,  tpd_A_SIGNEXTOUT(5), true),
						6 => (A_ipd(6)'last_event,  tpd_A_SIGNEXTOUT(6), true),
						7 => (A_ipd(7)'last_event,  tpd_A_SIGNEXTOUT(7), true),
						8=> (A_ipd(8)'last_event,  tpd_A_SIGNEXTOUT(8 ), true),
						9 => (A_ipd(9)'last_event,  tpd_A_SIGNEXTOUT(9), true),
						10 => (A_ipd(10)'last_event,  tpd_A_SIGNEXTOUT(10 ), true),
						11 => (A_ipd(11)'last_event,  tpd_A_SIGNEXTOUT(11), true),
						12 => (A_ipd(12)'last_event,  tpd_A_SIGNEXTOUT(12 ), true),
						13=> (A_ipd(13)'last_event,  tpd_A_SIGNEXTOUT(13), true),
						14=> (A_ipd(14)'last_event,  tpd_A_SIGNEXTOUT(14), true), 
						15=> (A_ipd(15)'last_event,  tpd_A_SIGNEXTOUT(15 ), true)
						),
      Mode          => VitalTransport,					
	  IgnoreDefaultDelay => TRUE,						  
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning); 
	  
	  
	  	   VitalPathDelay01 (
      OutSignal     => SIGNEXTOUT,
      GlitchData    => SIGNEXTOUT_GlitchData,
      OutSignalName => "SIGNEXTOUT",
      OutTemp       => SIGNEXTOUT_zd,
      Paths         => (0 => (B_ipd(0)'last_event,  tpd_B_SIGNEXTOUT(0), true),
						1 => (B_ipd(1)'last_event,  tpd_B_SIGNEXTOUT(1), true),
						2 => (B_ipd(2)'last_event,  tpd_B_SIGNEXTOUT(2), true),
						3 => (B_ipd(3)'last_event,  tpd_B_SIGNEXTOUT(3), true),
						4 => (B_ipd(4)'last_event,  tpd_B_SIGNEXTOUT(4), true), 
						5 => (B_ipd(5)'last_event,  tpd_B_SIGNEXTOUT(5), true),
						6 => (B_ipd(6)'last_event,  tpd_B_SIGNEXTOUT(6), true),
						7 => (B_ipd(7)'last_event,  tpd_B_SIGNEXTOUT(7), true),
						8=> (B_ipd(8)'last_event,  tpd_B_SIGNEXTOUT(8 ), true),
						9 => (B_ipd(9)'last_event,  tpd_B_SIGNEXTOUT(9), true),
						10 => (B_ipd(10)'last_event,  tpd_B_SIGNEXTOUT(10 ), true),
						11 => (B_ipd(11)'last_event,  tpd_B_SIGNEXTOUT(11), true),
						12 => (B_ipd(12)'last_event,  tpd_B_SIGNEXTOUT(12 ), true),
						13=> (B_ipd(13)'last_event,  tpd_B_SIGNEXTOUT(13), true),
						14=> (B_ipd(14)'last_event,  tpd_B_SIGNEXTOUT(14), true), 
						15=> (B_ipd(15)'last_event,  tpd_B_SIGNEXTOUT(15 ), true)
						),
      Mode          => VitalTransport,					
	  IgnoreDefaultDelay => TRUE,						  
	  RejectFastPath=>TRUE,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning); 
	  
	  
	end process VITALPathDelay;	

	mac16physical_i : mac16_physical  port map (
	 	CLK 	=> CLK_ipd,
	 	A	=> A_ipd,
	 	B	=> B_ipd,
	 	C	=> C_ipd,
	 	D	=> D_ipd,
	 	IHRST 	=> IRSTTOP_ipd,
	 	ILRST	=> IRSTBOT_ipd,
	 	OHRST	=> ORSTTOP_ipd,
	 	OLRST	=> ORSTBOT_ipd,
	 	AHLD	=> AHOLD_ipd,
	 	BHLD	=> BHOLD_ipd,
	 	CHLD	=> CHOLD_ipd,
	 	DHLD	=> DHOLD_ipd,		
	 	OHHLD	=> OHOLDTOP_ipd,
	 	OLHLD	=> OHOLDBOT_ipd,
	 	OHADS	=> ADDSUBTOP_ipd,
	 	OLADS	=> ADDSUBBOT_ipd,
	 	OHLDA	=> OLOADTOP_ipd,
	 	OLLDA	=> OLOADBOT_ipd,
	 	CICAS	=> ACCUMCI_ipd,
	 	CI		=> CI_ipd,
	 	SIGNEXTIN	=> SIGNEXTIN_ipd,
	 	SIGNEXTOUT	=> SIGNEXTOUT_zd,
	 	COCAS		=> QACCUMCO_zd,
	 	CO			=> QCO_zd,
	 	O			=> Q_zd , 
	 	CBIT		=> cbitss
    );

end  SB_MAC16_V; --SB_MAC16 


----------------------------------------------------------------
--		-- SB_IO_DLY --				     --- 
----------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all; 
use work.std_logic_SBT.all;
 
entity SB_IO_DLY is
	generic	(

		NEG_TRIGGER 		: bit				:='0';
		PIN_TYPE		: bit_vector (5 downto 0)	:="000000";
		PULLUP			: bit				:='0';
		IO_STANDARD		: string			:="SB_LVCMOS";
		INDELAY_VAL		: bit_vector (5 downto 0) 	:="000000";
		OUTDELAY_VAL 		: bit_vector (5 downto 0) 	:="000000"
	);	
	port 	(
		PACKAGE_PIN 		: inout std_ulogic; 
		LATCH_INPUT_VALUE 	: in 	std_logic; 
		CLOCK_ENABLE		: in 	std_logic; 
		INPUT_CLK		: in 	std_logic; 
		OUTPUT_CLK		: in 	std_logic; 
		OUTPUT_ENABLE		: in 	std_logic :='H'; 
		D_OUT_1			: in 	std_logic;   
		D_OUT_0			: in 	std_logic;  
		D_IN_1			: out 	std_logic; 
		D_IN_0			: out 	std_logic; 
		SCLK			: in 	std_logic; 	
		SDI			: in 	std_logic; 	
		C_R_SEL			: in 	std_logic;  
		SDO			: out 	std_logic 
	 );


end SB_IO_DLY; 	--  SB_IO_DLY 


architecture SB_IO_DLY_V of SB_IO_DLY is

	component	preio_physical
	port	(
			hold	:	in 	std_logic;
			rstio	:	in	std_logic;
			bs_en	:	in	std_logic;
			shift	:	in	std_logic;
			tclk	:	in	std_logic;
			inclk	:	in	std_logic;
			outclk	:	in	std_logic;
			update	:	in	std_logic;
			oepin	:	in	std_logic;
			sdi		:	in	std_logic;
			mode	:	in	std_logic;
			hiz_b	:	in	std_logic;
			sdo		:	out	std_logic;
			dout1	:	out	std_logic;
			dout0	:	out	std_logic;
			ddr1	:	in	std_logic;
			ddr0	:	in	std_logic;
			padin	:	in	std_logic;
			padout	:	out	std_logic;
			padoen	:	out	std_logic;
			cbit	:	in	std_logic_vector	(5 downto 0)
			);
	end component;	   
	
	component inoutdly64  
	generic ( 
		 INDELAY  		: bit_vector(5 downto 0)	:="000000"; 
		 OUTDELAY 		: bit_vector(5 downto 0) 	:="000000"  		 
	);
	port (
		sclk			: in 	std_logic := 'X';
		serialreg_rst   	: in  	std_logic := '1'; 				 
		sdi 			: in    std_logic := 'X';
		c_r_sel 		: in	std_logic := 'X';
		in_datain 		: in 	std_logic;
		out_datain 		: in  	std_logic;
		delay_direction		: in 	std_logic ; 
		delayed_dataout 	: out 	std_logic ; 
		sdo			: out 	std_logic := 'Z' 
	); 
	end component; 	
	
	signal	inclk_n, outclk_n, inclk, outclk,sdo_preio	:	std_logic;
	
	signal	bs_en	:	std_logic	:='0';	--Boundary scan enable           
	signal	shift	:	std_logic	:='0';	--Boundary scan shift            
	signal	tclk	:	std_logic	:='0';	--Boundary scan clock            
	signal	update	:	std_logic	:='0';	--Boundary scan update           
	signal	sdi_preio		:	std_logic	:='0';	--Boundary scan serial data in   
	signal	mode	:	std_logic	:='0';	--Boundary scan mode             
	signal	hiz_b	:	std_logic	:='1';	--Boundary scan Tristate control 
	
	signal	pin_cbit:	std_logic_vector(5 downto 0);
	signal	neg_trig:	std_logic;
	signal	pull_up	:	std_logic;
	signal	hold,oepin,padoen,padout,padin	:	std_logic;
	signal 	padinout_delayed 		: 	std_logic; 
	signal  INCLKE_sync , OUTCLKE_sync     : std_logic; 
begin
	
	pin_cbit	<=	TO_STDLOGICVECTOR	(PIN_TYPE);
	neg_trig	<=	TO_STDLOGIC	(NEG_TRIGGER);
	pull_up		<=	TO_STDLOGIC	(PULLUP);

	inclk_n	<= 	INPUT_CLK xor neg_trig;
	outclk_n<=	OUTPUT_CLK xor neg_trig;
--	inclk	<=	inclk_n and CLOCK_ENABLE;
--	outclk	<=	outclk_n and CLOCK_ENABLE;

	process(inclk_n , CLOCK_ENABLE) is         begin
                if(inclk_n ='0') then
                        INCLKE_sync  <= CLOCK_ENABLE;
                else
                        INCLKE_sync <= INCLKE_sync;
                end if ;
        end process;

        process(outclk_n , CLOCK_ENABLE) is
        begin
                if(outclk_n ='0') then
                        OUTCLKE_sync  <= CLOCK_ENABLE;
                else
                        OUTCLKE_sync <= OUTCLKE_sync;
                end if ;
        end process;

        inclk <= (inclk_n and INCLKE_sync);
        outclk <= (outclk_n and OUTCLKE_sync);

	
	hold	<=	LATCH_INPUT_VALUE;
	oepin	<=	OUTPUT_ENABLE;
	
	PACKAGE_PIN_i	:	process	(padoen, padinout_delayed, PACKAGE_PIN)
	begin
		padin	<=	PACKAGE_PIN;
		if	(padoen='1') then
			PACKAGE_PIN	<=	'Z';
		else
			PACKAGE_PIN	<=	padinout_delayed;
		end if;
	end process;
-----------------------------------------------------------------	
	preio_physical_i	:	preio_physical
	port map	(
				hold	=>	hold,
				rstio	=>	'0',
				bs_en	=>	bs_en,
				shift	=>	shift,
				tclk	=>	tclk,
				inclk	=>	inclk,
				outclk	=>	outclk,
				update	=>	update,
				oepin	=>	oepin,
				sdi		=>	sdi_preio,
				mode	=>	mode,
				hiz_b	=>	hiz_b,
				sdo		=>	sdo_preio,
				dout1	=>	D_IN_1,
				dout0	=>	D_IN_0,
				ddr1	=>	D_OUT_1,
				ddr0	=>	D_OUT_0,
				padin	=>	padinout_delayed,
				padout	=>	padout,
				padoen	=>	padoen,
				cbit	=>	pin_cbit
				);
				
	inoutdly64_i  : inoutdly64 
	generic map  ( 
		 INDELAY  		=> INDELAY_VAL ,  
		 OUTDELAY 		=> OUTDELAY_VAL
	)
	port map (
		-- disabled dynamic delay test logic sections
		sclk			=>open,
		serialreg_rst   	=>open, 
		sdi 			=>open,  
		c_r_sel 		=>open, 
		in_datain 		=> padin,
		out_datain 		=> padout, 
		delay_direction		=> padoen,   
		delayed_dataout 	=> padinout_delayed, 
		sdo			=> open); 
	
end SB_IO_DLY_V;

---------------------------------------------------------------------------
----			 	inoutdly64  				---	
---------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;
 

entity inoutdly64  is
 
	generic ( 
		 INDELAY  			: bit_vector(5 downto 0)	:="000000"; 
		 OUTDELAY 			: bit_vector(5 downto 0) 	:="000000"  		 
	);
	port (
		sclk		: in 	std_logic;
		serialreg_rst   : in  	std_logic; 				 
		sdi 		: in    std_logic; 
		c_r_sel 	: in	std_logic;
		in_datain 	: in 	std_logic;
		out_datain 	: in  	std_logic;
		delay_direction	: in 	std_logic ; 
		delayed_dataout : out 	std_logic ; 
		sdo		: out 	std_logic 
	); 

end inoutdly64;
	
architecture inoutdly64_arch  of inoutdly64 is

-- signal for generics  
signal	indelay_generic 			: std_logic_vector( 5 downto 0);  
signal	outdelay_generic  			: std_logic_vector( 5 downto 0);  
-- logic signals 
signal  serial_data				: std_logic_vector(11 downto 0):="000000000000";
signal  buf_y					: std_logic_vector(63 downto 0) ; 
signal  data_in 				: std_logic; 
signal  delayval_sel				: std_logic_vector(5 downto 0); 
signal  delayed_data				: std_logic;   

begin 
	-- generic to signal conversions --  	
	indelay_generic 		<= TO_STDLOGICVECTOR(INDELAY); 
	outdelay_generic 		<= TO_STDLOGICVECTOR(OUTDELAY);				

	-- logic section ---  		
	serialdata_proc:  process (sclk,serialreg_rst) is 
		begin 
		if(serialreg_rst = '1') then 	 
			serial_data <= (Others  => '0'); 
		elsif rising_edge(sclk) then
			serial_data <= sdi & serial_data(11 downto 1);
		end if;
	end process;

	sdo <= serial_data(0); 	 	
			
	seldatain_proc : process(delay_direction, in_datain,out_datain) 
		begin 
		case delay_direction is 
		when '0' => data_in <= out_datain ;  -- preio_oen =0
		when '1' => data_in <= in_datain ;   -- preio_oen =1 
		when others => data_in <= out_datain ;
		end case;  
	end process; 	

	-- dynamic delay selection & shiftreg delay logics are not required. Static delays are applied through in,out parameters 
	--seldelaytype_proc: process(delay_direction, c_r_sel,indelay_generic, outdelay_generic,serial_data) 
	--	variable seldelaydata :  std_logic_vector( 1 downto 0); 
	--	begin 
	--	seldelaydata :=(delay_direction & c_r_sel);
	--	case seldelaydata is 
	--		when "00" => 
	--			delayval_sel <= outdelay_generic(5 downto 0);		-- out line delay static 
	--		when "01" => 
	--			delayval_sel <= serial_data(11 downto 6);       -- out line delay dynamic 
	--		when "10" => 
	--			delayval_sel <= indelay_generic(5 downto 0);     -- in line delay static 
	--		when "11" => 
	--			delayval_sel <= serial_data(5 downto 0);        -- in line delay dynamic 
	--		when others =>
	--			delayval_sel <= (others => '0');         
	--		end case ; 
	--end process; 

	-- Static delay selection 
	seldelayval_static_proc : process(delay_direction, indelay_generic, outdelay_generic)  
		begin 
		case delay_direction is 
		when '0' => delayval_sel  <= outdelay_generic ;  -- preio_oen =0
		when '1' => delayval_sel  <= indelay_generic  ;   -- preio_oen =1 
		when others => delayval_sel  <= outdelay_generic ;
		end case;  
	end process; 	

	-- delay tap  generation  	
	buf_y(0) <= data_in; 	
	delaytap_gen: for N in 1 to 63 generate 
	buf_y(N) <= buf_y(N-1) after  100 ps ;             -- 100ps +-25ps.  
	end generate;

	seldelayeddata_proc: process(delayval_sel,buf_y ) 
	begin				  
		delayed_data <=buf_y(slv_to_integer(delayval_sel)); 
	end process;   
	
	delayed_dataout <= delayed_data; 	
 
end inoutdly64_arch;

------------------------------------------------------------------
--	 SB_MIPI_TX_4LANE				      	--
------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;
 
entity SB_MIPI_TX_4LANE is

	generic	( 		
		DIVR 			: bit_vector( 4 downto 0)  	:= "11111" ;      	-- Ref Clk divider
		DIVF 			: bit_vector( 7 downto 0)  	:= "11110000"; 		-- Feedback divider
		DIVQ 			: bit_vector( 1 downto 0)  	:= "00";       		-- VCO divider
		TEST_MODE 		: bit 				:= '0';
		TEST_BITS 		: bit_vector( 3 downto 0) 	:= "1001"
	); 
	port 	( 
			--Common Interface Pins
		PU			: in 	std_logic ; 
		LBEN			: in 	std_logic ; 
 		ROUTCAL			: in 	std_logic_vector(1 downto 0) ; 
 		ENPDESER		: in	std_logic ; 	
	       	PDCKG			: in	std_logic ; 
			-- DATA0 Interface pins
		DP0			: inout	std_ulogic ; 	
		DN0			: inout std_ulogic ; 
 		D0OPMODE		: in	std_logic ;  
 		D0DTXLPP		: in	std_logic ; 
 		D0DTXLPN		: in 	std_logic ; 
 		D0TXLPEN		: in	std_logic ;  	
 		D0DRXLPP		: out	std_logic ; 
	  	D0DRXLPN		: out 	std_logic ; 
 		D0RXLPEN		: in 	std_logic ; 
 		D0DCDP			: out 	std_logic ; 
		D0DCDN			: out 	std_logic ; 
 		D0CDEN			: in	std_logic ; 		
  		D0TXHSPD		: in	std_logic ; 
 		D0TXHSEN		: in 	std_logic ; 
   		D0HSTXDATA		: in 	std_logic_vector( 7 downto 0) ; 
  		D0HSSEREN		: in	std_logic ; 	 
 		D0RXHSEN		: in	std_logic ; 
  		D0HSDESEREN		: in 	std_logic ; 	
 	 	D0HSRXDATA		: out 	std_logic_vector( 7 downto 0) ; 
 		D0HSBYTECLKD		: out 	std_logic ; 
 		D0SYNC			: out 	std_logic ; 
 		D0ERRSYNC		: out 	std_logic ; 
	      	D0HSBYTECLKSNOSYNC	: out 	std_logic ; 
			-- DATA1 Interface pins
		DP1			: inout std_ulogic ; 
		DN1			: inout std_ulogic ;  
 		D1DTXLPP		: in 	std_logic ; 
 		D1DTXLPN		: in	std_logic ; 
  		D1TXLPEN		: in 	std_logic ; 
 		D1DRXLPP		: out 	std_logic ;
	  	D1DRXLPN		: out 	std_logic ; 
 		D1RXLPEN		: in	std_logic ;
 		D1DCDP			: out 	std_logic ; 
		D1DCDN			: out  	std_logic ; 
 		D1CDEN			: in	std_logic ; 
  		D1TXHSPD		: in 	std_logic ; 
 		D1TXHSEN		: in	std_logic ;  
		D1HSTXDATA		: in 	std_logic_vector( 7 downto 0) ; 
  		D1HSSEREN		: in	std_logic ; 
 		D1RXHSEN		: in 	std_logic ;
  		D1HSDESEREN		: in 	std_logic ; 
	 	D1HSRXDATA		: out   std_logic_vector( 7 downto 0) ; 
 		D1SYNC			: out 	std_logic ; 
 		D1ERRSYNC		: out 	std_logic ; 
 		D1NOSYNC		: out 	std_logic ; 
			-- DATA2 Interface pins
		DP2			: inout std_ulogic ;
		DN2			: inout std_ulogic ; 
 		D2DTXLPP		: in	std_logic ; 
 		D2DTXLPN		: in 	std_logic ; 
  		D2TXLPEN		: in 	std_logic ; 
 		D2DRXLPP		: out 	std_logic ; 
	  	D2DRXLPN		: out 	std_logic ; 
 		D2RXLPEN		: in 	std_logic ; 
 		D2DCDP			: out 	std_logic ; 
		D2DCDN			: out 	std_logic ; 
 		D2CDEN			: in	std_logic ;
  		D2TXHSPD		: in	std_logic ; 
 		D2TXHSEN		: in	std_logic ; 		 
    	 	D2HSTXDATA		: in	std_logic_vector( 7 downto 0) ; 
  		D2HSSEREN		: in	std_logic ; 
 		D2RXHSEN		: in	std_logic ; 
  		D2HSDESEREN		: in	std_logic ; 
 	 	D2HSRXDATA		: out 	std_logic_vector( 7 downto 0) ; 
 		D2SYNC			: out 	std_logic ; 
 		D2ERRSYNC		: out 	std_logic ;
 		D2NOSYNC		: out 	std_logic ; 
			-- DATA3 Interface pins
		DP3			: inout std_ulogic ; 
		DN3			: inout std_ulogic ;
 		D3DTXLPP		: in 	std_logic ; 
 		D3DTXLPN		: in	std_logic ; 
  		D3TXLPEN		: in 	std_logic ; 
 		D3DRXLPP		: out 	std_logic ; 
	  	D3DRXLPN		: out 	std_logic ;
 		D3RXLPEN		: in	std_logic ; 
 		D3DCDP			: out 	std_logic ; 
		D3DCDN			: out 	std_logic ; 
 		D3CDEN			: in	std_logic ; 
  		D3TXHSPD		: in	std_logic ; 
 		D3TXHSEN		: in	std_logic ;  
  	 	D3HSTXDATA		: in 	std_logic_vector( 7 downto 0) ; 
  		D3HSSEREN		: in	std_logic ; 
 		D3RXHSEN		: in	std_logic ; 
  		D3HSDESEREN		: in	std_logic ; 
 	 	D3HSRXDATA		: out 	std_logic_vector( 7 downto 0) ; 
 		D3SYNC			: out 	std_logic ;	
 		D3ERRSYNC		: out	std_logic ; 
 		D3NOSYNC		: out 	std_logic ; 
			-- CLOCK Interface pins
		CKP			: inout std_ulogic ;  	
		CKN			: inout std_ulogic ;   
 		CLKDTXLPP		: in 	std_logic ; 
 		CLKDTXLPN		: in	std_logic ; 
  		CLKTXLPEN		: in 	std_logic ; 
	  	CLKDRXLPP		: out 	std_logic ; 
	  	CLKDRXLPN		: out 	std_logic ; 
  		CLKRXLPEN		: in	std_logic ; 
  		CLKTXHSPD		: in	std_logic ; 
 		CLKTXHSEN		: in	std_logic ; 
	       	CLKTXHSGATE		: in	std_logic ; 
  		CLKRXHSEN		: in	std_logic ; 
	     	CLKHSBYTE		: out 	std_logic ; 
			-- Universal MIPI PLL Interface pins
 		PLLPU			: in 	std_logic ; 
 		PLLREF			: in	std_logic ; 
 		PLLLOCK			: out 	std_logic ; 
			-- Universal MIPI PLL Serial Configuration Register Interface pins
 		PLLCFGSRDI		: in	std_logic ; 
 		PLLCFGSRRESET		: in	std_logic ; 
 		PLLCFGSRCLK		: in	std_logic ; 
 		PLLCFGSRDO		: out 	std_logic 
	);

	-- Device Pins: DP3,DN3,DP2,DN2,DP1,DN1,DP0,DN0,CKP,CKN.

end SB_MIPI_TX_4LANE;  -- SB_MIPI_TX_4LANE 

architecture SB_MIPI_TX_4LANE_V  of SB_MIPI_TX_4LANE  is

component  X1082T001 is 
port (
		---- Power Pins 
        	VDDA 		: in		std_logic;
           	VSSA		: in		std_logic;
	        VDD		: in 		std_logic;
        	VSS		: in		std_logic;
	        DVSS		: in		std_logic;
		---- Common Interface Pins
	        BITCLK		: in 		std_logic;
 		PD		: in 		std_logic;
		LB_EN		: in		std_logic;
 		ROUT_CAL	: in 		std_logic_vector(1 downto 0);
 		ENP_DESER	: in		std_logic;
           	PDCKG		: in		std_logic;
		----  DATA0 Interface pins
  		DP0		: inout 	std_logic ; 
	  	DN0		: inout 	std_logic ;
		D0_OPMODE	: in		std_logic ;
		D0_DTXLPP	: in		std_logic ;
		D0_DTXLPN	: in		std_logic ;
 		D0_TXLPEN	: in 		std_logic ;
 		D0_DRXLPP	: out		std_logic ;
	  	D0_DRXLPN	: out		std_logic ;
		D0_RXLPEN	: in		std_logic ;
 		D0_DCDP		: out 		std_logic ;
		D0_DCDN		: out           std_logic ;
		D0_CDEN		: in    	std_logic ;
 		D0_TXHSPD	: in    	std_logic ;
		D0_TXHSEN	: in    	std_logic ;
		D0_HSTX_DATA	: in    	std_logic_vector(7 downto 0) ;
 		D0_HS_SER_EN	: in    	std_logic ;
		D0_RXHSEN	: in    	std_logic ;
 		D0_HS_DESER_EN	: in    	std_logic ;
 	 	D0_HSRX_DATA 	: out           std_logic_vector( 7 downto 0);
 		D0_HS_BYTE_CLKD : out           std_logic ;
 		D0_SYNC		: out           std_logic ;
 		D0_ERRSYNC	: out           std_logic ;
         	D0_HS_BYTE_CLKS_NOSYNC	: out 	std_logic ;
		----  DATA1 Interface pins
	  	DP1		: inout    	std_logic;
  		DN1		: inout    	std_logic;
		D1_DTXLPP	: in    	std_logic;
		D1_DTXLPN	: in    	std_logic;
 		D1_TXLPEN	: in    	std_logic;
 		D1_DRXLPP	: out    	std_logic;
	  	D1_DRXLPN	: out    	std_logic;
		D1_RXLPEN	: in    	std_logic;
 		D1_DCDP		: out    	std_logic;
		D1_DCDN		: out    	std_logic;
		D1_CDEN		: in    	std_logic;
 		D1_TXHSPD	: in    	std_logic;
		D1_TXHSEN	: in    	std_logic; 
   	 	D1_HSTX_DATA	: in    	std_logic_vector(7 downto 0);
 		D1_HS_SER_EN	: in    	std_logic;
		D1_RXHSEN	: in    	std_logic;
 		D1_HS_DESER_EN	: in    	std_logic;
 	 	D1_HSRX_DATA	: out    	std_logic_vector(7 downto 0);
 		D1_SYNC		: out    	std_logic;
 		D1_ERRSYNC	: out    	std_logic;
 		D1_NOSYNC 	: out    	std_logic;
		----  DATA2 Interface pins
	  	DP2 		: inout    	std_logic ;
  		DN2 		: inout    	std_logic ;
		D2_DTXLPP	: in    	std_logic ;
		D2_DTXLPN	: in    	std_logic ;
 		D2_TXLPEN	: in    	std_logic ;
 		D2_DRXLPP	: out    	std_logic ;
	  	D2_DRXLPN	: out    	std_logic ;
		D2_RXLPEN 	: in    	std_logic ;
 		D2_DCDP	 	: out    	std_logic ;
		D2_DCDN 	: out    	std_logic ;
		D2_CDEN 	: in    	std_logic ;
 		D2_TXHSPD 	: in    	std_logic ;
		D2_TXHSEN 	: in    	std_logic ; 
   		D2_HSTX_DATA 	: in    	std_logic_vector(7 downto 0) ;
 		D2_HS_SER_EN 	: in    	std_logic ;
		D2_RXHSEN 	: in    	std_logic ;
 		D2_HS_DESER_EN 	: in    	std_logic ;
 	 	D2_HSRX_DATA 	: out    	std_logic_vector(7 downto 0);
 		D2_SYNC 	: out   	std_logic;
 		D2_ERRSYNC 	: out    	std_logic;
 		D2_NOSYNC 	: out    	std_logic ;
		---- DATA3 Interface pins
	  	DP3 		: inout    	std_logic;
  		DN3 		: inout    	std_logic;
		D3_DTXLPP 	: in    	std_logic;
		D3_DTXLPN 	: in    	std_logic;
 		D3_TXLPEN 	: in    	std_logic ;
 		D3_DRXLPP 	: out    	std_logic;
	  	D3_DRXLPN 	: out    	std_logic ;
		D3_RXLPEN 	: in    	std_logic;
 		D3_DCDP 	: out    	std_logic;
		D3_DCDN 	: out    	std_logic;
		D3_CDEN 	: in    	std_logic;
 		D3_TXHSPD 	: in    	std_logic ;
		D3_TXHSEN 	: in    	std_logic; 
   		D3_HSTX_DATA 	: in    	std_logic_vector(7 downto 0);
 		D3_HS_SER_EN 	: in    	std_logic;
		D3_RXHSEN 	: in    	std_logic ;
 		D3_HS_DESER_EN 	: in    	std_logic ;
 	 	D3_HSRX_DATA 	: out    	std_logic_vector(7 downto 0);
 		D3_SYNC 	: out    	std_logic ;
 		D3_ERRSYNC 	: out    	std_logic ;
 		D3_NOSYNC 	: out    	std_logic ;
		---- CLOCK Interface pins
	  	CKP 		: inout 	std_logic ;
  		CKN 		: inout  	std_logic ;
		CLK_DTXLPP 	: in   	 	std_logic ;
		CLK_DTXLPN 	: in    	std_logic ;
 		CLK_TXLPEN 	: in   	 	std_logic ;
	  	CLK_DRXLPP 	: out    	std_logic ;
  		CLK_DRXLPN 	: out    	std_logic ;
 		CLK_RXLPEN 	: in    	std_logic ;
 		CLK_TXHSPD 	: in    	std_logic ;
		CLK_TXHSEN 	: in    	std_logic ;
	        CLK_TXHSGATE 	: in    	std_logic ;
 		CLK_RXHSEN 	: in   	 	std_logic ;
        	CLK_HS_BYTE 	: out    	std_logic 
		); 
end component; 

component  X109T001 is  
port ( 
		VDDA		: in		std_logic ; 
		VSSA		: in            std_logic ;
		VDD 		: in            std_logic ;
		VSS		: in            std_logic ;
		PD		: in            std_logic ;	       			--  Power Down, active high
		TST	 	: in            std_logic_vector(3 downto 0) ;		
		CN		: in            std_logic_vector(4 downto 0) ;		--  Control N divider
		CM		: in            std_logic_vector(7 downto 0) ;		--  Control M divider
		CO		: in            std_logic_vector(1 downto 0) ;		--  Control O divider
		CLKREF	        : in            std_logic ;				--  Reference clock input
		OUTP	        : out           std_logic ;				--  Output clock (P)
		OUTN	        : out           std_logic ;				--  Output clock (N)
		LOCK	        : out 	 	std_logic 				--   Lock detection. When high, the PLL has achieved
); 
end component; 

	signal divr_gen 	: std_logic_vector( 4 downto 0);
	signal divf_gen 	: std_logic_vector( 7 downto 0); 
	signal divq_gen 	: std_logic_vector( 1 downto 0); 
	signal testmode 	: std_logic; 
	signal testbits 	: std_logic_vector( 3 downto 0);  

	signal BITCLK_int 	: std_logic;
	signal not_PU 		: std_logic;  
	signal not_PLLPU	: std_logic; 

begin 
	-- generic to signal conversion 
	divr_gen	<= TO_STDLOGICVECTOR(DIVR);   
	divf_gen 	<= TO_STDLOGICVECTOR(DIVF); 
	divq_gen  	<= TO_STDLOGICVECTOR(DIVQ); 
	testmode	<= TO_STDLOGIC(TEST_MODE); 	
 	testbits 	<= TO_STDLOGICVECTOR(TEST_BITS); 

	not_PU <= not(PU); 
	not_PLLPU <= not(PLLPU); 

	mipi_txrxphy_i 		:   X1082T001  
	port map  (
		---- Power Pins 
        	VDDA 		=> '1' ,
           	VSSA		=> '0' ,
	        VDD		=> '1' ,
        	VSS		=> '0' , 
	        DVSS		=> '0' , 
		---- Common Interface Pins
	        BITCLK		=> BITCLK_int , 
 		PD		=> not_PU,  
		LB_EN		=> LBEN ,
 		ROUT_CAL	=> ROUTCAL ,
 		ENP_DESER	=> ENPDESER ,
           	PDCKG		=> PDCKG ,
		----  DATA0 Interface pins
  		DP0		=> DP0 , 
	  	DN0		=> DN0 ,
		D0_OPMODE	=> D0OPMODE ,
		D0_DTXLPP	=> D0DTXLPP ,
		D0_DTXLPN	=> D0DTXLPN ,
 		D0_TXLPEN	=> D0TXLPEN ,
 		D0_DRXLPP	=> D0DRXLPP ,
	  	D0_DRXLPN	=> D0DRXLPN ,
		D0_RXLPEN	=> D0RXLPEN ,
 		D0_DCDP		=> D0DCDP ,
		D0_DCDN		=> D0DCDN ,
		D0_CDEN		=> D0CDEN ,
 		D0_TXHSPD	=> D0TXHSPD ,
		D0_TXHSEN	=> D0TXHSEN  ,
		D0_HSTX_DATA	=> D0HSTXDATA ,
 		D0_HS_SER_EN	=> D0HSSEREN ,
		D0_RXHSEN	=> D0RXHSEN ,
 		D0_HS_DESER_EN	=> D0HSDESEREN ,
 	 	D0_HSRX_DATA 	=> D0HSRXDATA ,
 		D0_HS_BYTE_CLKD => D0HSBYTECLKD ,
 		D0_SYNC		=> D0SYNC ,
 		D0_ERRSYNC	=> D0ERRSYNC ,
         	D0_HS_BYTE_CLKS_NOSYNC	=> D0HSBYTECLKSNOSYNC ,
		----  DATA1 Interface pins
	  	DP1		=> DP1 ,
  		DN1		=> DN1 ,
		D1_DTXLPP	=> D1DTXLPP ,
		D1_DTXLPN	=> D1DTXLPN ,
 		D1_TXLPEN	=> D1TXLPEN ,
 		D1_DRXLPP	=> D1DRXLPP ,
	  	D1_DRXLPN	=> D1DRXLPN ,
		D1_RXLPEN	=> D1RXLPEN ,
 		D1_DCDP		=> D1DCDP ,
		D1_DCDN		=> D1DCDN ,
		D1_CDEN		=> D1CDEN ,
 		D1_TXHSPD	=> D1TXHSPD ,
		D1_TXHSEN	=> D1TXHSEN , 
   	 	D1_HSTX_DATA	=> D1HSTXDATA ,
 		D1_HS_SER_EN	=> D1HSSEREN ,
		D1_RXHSEN	=> D1RXHSEN ,
 		D1_HS_DESER_EN	=> D1HSDESEREN ,
 	 	D1_HSRX_DATA	=> D1HSRXDATA ,
 		D1_SYNC		=> D1SYNC ,
 		D1_ERRSYNC	=> D1ERRSYNC ,
 		D1_NOSYNC 	=> D1NOSYNC ,
		----  DATA2 Interface pins
	  	DP2 		=> DP2 ,
  		DN2 		=> DN2 ,
		D2_DTXLPP	=> D2DTXLPP ,
		D2_DTXLPN	=> D2DTXLPN ,
 		D2_TXLPEN	=> D2TXLPEN ,
 		D2_DRXLPP	=> D2DRXLPP ,
	  	D2_DRXLPN	=> D2DRXLPN ,
		D2_RXLPEN 	=> D2RXLPEN ,
 		D2_DCDP	 	=> D2DCDP ,
		D2_DCDN 	=> D2DCDN ,
		D2_CDEN 	=> D2CDEN ,
 		D2_TXHSPD 	=> D2TXHSPD ,
		D2_TXHSEN 	=> D2TXHSEN , 
   		D2_HSTX_DATA 	=> D2HSTXDATA ,
 		D2_HS_SER_EN 	=> D2HSSEREN ,
		D2_RXHSEN 	=> D2RXHSEN  ,
 		D2_HS_DESER_EN 	=> D2HSDESEREN ,
 	 	D2_HSRX_DATA 	=> D2HSRXDATA ,
 		D2_SYNC 	=> D2SYNC ,
 		D2_ERRSYNC 	=> D2ERRSYNC ,
 		D2_NOSYNC 	=> D2NOSYNC ,
		---- DATA3 Interface pins
	  	DP3 		=> DP3 ,
  		DN3 		=> DN3 ,
		D3_DTXLPP 	=> D3DTXLPP ,
		D3_DTXLPN 	=> D3DTXLPN ,
 		D3_TXLPEN 	=> D3TXLPEN ,
 		D3_DRXLPP 	=> D3DRXLPP ,
	  	D3_DRXLPN 	=> D3DRXLPN ,
		D3_RXLPEN 	=> D3RXLPEN ,
 		D3_DCDP 	=> D3DCDP ,
		D3_DCDN 	=> D3DCDN ,
		D3_CDEN 	=> D3CDEN ,
 		D3_TXHSPD 	=> D3TXHSPD ,
		D3_TXHSEN 	=> D3TXHSEN , 
   		D3_HSTX_DATA 	=> D3HSTXDATA ,
 		D3_HS_SER_EN 	=> D3HSSEREN ,
		D3_RXHSEN 	=> D3RXHSEN ,
 		D3_HS_DESER_EN 	=> D3HSDESEREN ,
 	 	D3_HSRX_DATA 	=> D3HSRXDATA ,
 		D3_SYNC 	=> D3SYNC ,
 		D3_ERRSYNC 	=> D3ERRSYNC ,
 		D3_NOSYNC 	=> D3NOSYNC ,
		---- CLOCK Interface pins
	  	CKP 		=> CKP ,
  		CKN 		=> CKN ,
		CLK_DTXLPP 	=> CLKDTXLPP  ,
		CLK_DTXLPN 	=> CLKDTXLPN  ,
 		CLK_TXLPEN 	=> CLKTXLPEN  ,
	  	CLK_DRXLPP 	=> CLKDRXLPP  ,
  		CLK_DRXLPN 	=> CLKDRXLPN  ,
 		CLK_RXLPEN 	=> CLKRXLPEN  ,
 		CLK_TXHSPD 	=> CLKTXHSPD  ,
		CLK_TXHSEN 	=> CLKTXHSEN  ,
	        CLK_TXHSGATE 	=> CLKTXHSGATE ,
 		CLK_RXHSEN 	=> CLKRXHSEN ,
        	CLK_HS_BYTE 	=> CLKHSBYTE  	 
		);

	
	mipi_txpllphy_i  : X109T001 
	port map (
		VDDA 		=> '1' ,
		VSSA 		=> '0' ,
		VDD 		=> '1' ,
		VSS 		=> '0' ,
		PD 		=> not_PLLPU , 
		TST 		=> "0000",        
		CN 		=> divr_gen,
		CM 		=> divf_gen,
		CO 		=> divq_gen,
		CLKREF 		=> PLLREF,
		OUTP 		=> BITCLK_int,
		OUTN 		=> open,
		LOCK 		=> PLLLOCK	
	 	);	
 

end SB_MIPI_TX_4LANE_V;

-----------------------------------------------------------------------------------------------------
--              	 ICE40MH 16K Block RAM Primitives  					   --  
-----------------------------------------------------------------------------------------------------
-- Front End Primitives :  
--	# SB_RAM1024x16		# SB_RAM1024x16NR  	# SB_RAM1024x16NW	# SB_RAM1024x16NRNW
--	# SB_RAM2048x8		# SB_RAM2048x8NR	# SB_RAM2048x8NW	# SB_RAM2048x8NRNW
--	# SB_RAM4096x4		# SB_RAM4096x4NR	# SB_RAM4096x4NW	# SB_RAM4096x4NRNW
--	# SB_RAM8192x2		# SB_RAM8192x2NR	# SB_RAM8192x2NW	# SB_RAM8192x2NRNW
-- Back End Primitives  : 
--	# SB_RAM40_16K		# SB_RAM40_16KNR 	# SB_RAM40_16KNW 	# SB_RAM40_16KNRNW
-------------------------------------------------------------------------------------------------------

---------------------------------------
	--- SB_RAM1024x16
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM1024x16 is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 
           INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 
           INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;

          port( 
                RDATA : out std_logic_vector( 15  downto 0) ;
                RCLK  : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'H';
                RADDR : in  std_logic_vector( 9  downto 0) ;
                WCLK  : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'H';
                WADDR : in  std_logic_vector( 9  downto 0) ;
                MASK  : in  std_logic_vector( 15  downto 0) ;
                WDATA : in  std_logic_vector( 15  downto 0)
               );
  
  
end SB_RAM1024x16;

architecture SB_RAM1024x16_ARCH of SB_RAM1024x16 is

  signal MEM : std_logic_vector(16383 downto 0) ;
  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLK)
  variable WADDR_in : integer range 0 to 1023;

    variable MEM_temp : std_logic_vector(16383 downto 0) :=  To_StdLogicVector(INIT_3F) &
                                                  To_StdLogicVector(INIT_3E) &
                                                  To_StdLogicVector(INIT_3D) &
                                                  To_StdLogicVector(INIT_3C) &
                                                  To_StdLogicVector(INIT_3B) &
                                                  To_StdLogicVector(INIT_3A) &
                                                  To_StdLogicVector(INIT_39) &
                                                  To_StdLogicVector(INIT_38) &
                                                  To_StdLogicVector(INIT_37) &
                                                  To_StdLogicVector(INIT_36) &
                                                  To_StdLogicVector(INIT_35) &
                                                  To_StdLogicVector(INIT_34) &
                                                  To_StdLogicVector(INIT_33) &
                                                  To_StdLogicVector(INIT_32) &
                                                  To_StdLogicVector(INIT_31) &
                                                  To_StdLogicVector(INIT_30) &
						  To_StdLogicVector(INIT_2F) &
                                                  To_StdLogicVector(INIT_2E) &
                                                  To_StdLogicVector(INIT_2D) &
                                                  To_StdLogicVector(INIT_2C) &
                                                  To_StdLogicVector(INIT_2B) &
                                                  To_StdLogicVector(INIT_2A) &
                                                  To_StdLogicVector(INIT_29) &
                                                  To_StdLogicVector(INIT_28) &
                                                  To_StdLogicVector(INIT_27) &
                                                  To_StdLogicVector(INIT_26) &
                                                  To_StdLogicVector(INIT_25) &
                                                  To_StdLogicVector(INIT_24) &
                                                  To_StdLogicVector(INIT_23) &
                                                  To_StdLogicVector(INIT_22) &
                                                  To_StdLogicVector(INIT_21) &
                                                  To_StdLogicVector(INIT_20) &
						  To_StdLogicVector(INIT_1F) &
                                                  To_StdLogicVector(INIT_1E) &
                                                  To_StdLogicVector(INIT_1D) &
                                                  To_StdLogicVector(INIT_1C) &
                                                  To_StdLogicVector(INIT_1B) &
                                                  To_StdLogicVector(INIT_1A) &
                                                  To_StdLogicVector(INIT_19) &
                                                  To_StdLogicVector(INIT_18) &
                                                  To_StdLogicVector(INIT_17) &
                                                  To_StdLogicVector(INIT_16) &
                                                  To_StdLogicVector(INIT_15) &
                                                  To_StdLogicVector(INIT_14) &
                                                  To_StdLogicVector(INIT_13) &
                                                  To_StdLogicVector(INIT_12) &
                                                  To_StdLogicVector(INIT_11) &
                                                  To_StdLogicVector(INIT_10) & 
						  To_StdLogicVector(INIT_F)  &
                                                  To_StdLogicVector(INIT_E)  &
                                                  To_StdLogicVector(INIT_D)  &
                                                  To_StdLogicVector(INIT_C)  &
                                                  To_StdLogicVector(INIT_B)  &
                                                  To_StdLogicVector(INIT_A)  &
                                                  To_StdLogicVector(INIT_9)  &
                                                  To_StdLogicVector(INIT_8)  &
                                                  To_StdLogicVector(INIT_7)  &
                                                  To_StdLogicVector(INIT_6)  &
                                                  To_StdLogicVector(INIT_5)  &
                                                  To_StdLogicVector(INIT_4)  &
                                                  To_StdLogicVector(INIT_3)  &
                                                  To_StdLogicVector(INIT_2)  &
                                                  To_StdLogicVector(INIT_1)  & 
                                                  To_StdLogicVector(INIT_0) ;  
  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLK'event and (WCLK = '1') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 15 loop
         if (MASK(i) = '0') then
            MEM_temp(16*WADDR_in + i )  := WDATA(i) ;
         end if ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;

  end process ;


  ReadBehavior : process(RCLK)
  
    variable RADDR_in : integer range 0 to 1023 ;
    variable RDATA_temp : std_logic_vector( 15  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLK'event and (RCLK = '1') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 15 loop
            RDATA_temp(i ) := MEM(16*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;

  end process ;

end SB_RAM1024x16_ARCH;   --- SB_RAM1024x16


---------------------------------------
	--- SB_RAM1024x16NR
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM1024x16NR is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 15  downto 0) ;
                RCLKN : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'H';
                RADDR : in  std_logic_vector( 9  downto 0) ;
                WCLK  : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'H';
                WADDR : in  std_logic_vector( 9  downto 0) ;
                MASK  : in  std_logic_vector( 15  downto 0) ;
                WDATA : in  std_logic_vector( 15  downto 0)
               );
  
  
end SB_RAM1024x16NR;

architecture SB_RAM1024x16NR_ARCH of SB_RAM1024x16NR is

  signal MEM : std_logic_vector(16383 downto 0) ;
  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLK)
  variable WADDR_in : integer range 0 to 1023;

    variable MEM_temp : std_logic_vector(16383 downto 0) :=  To_StdLogicVector(INIT_3F) &
                                                  To_StdLogicVector(INIT_3E) &
                                                  To_StdLogicVector(INIT_3D) &
                                                  To_StdLogicVector(INIT_3C) &
                                                  To_StdLogicVector(INIT_3B) &
                                                  To_StdLogicVector(INIT_3A) &
                                                  To_StdLogicVector(INIT_39) &
                                                  To_StdLogicVector(INIT_38) &
                                                  To_StdLogicVector(INIT_37) &
                                                  To_StdLogicVector(INIT_36) &
                                                  To_StdLogicVector(INIT_35) &
                                                  To_StdLogicVector(INIT_34) &
                                                  To_StdLogicVector(INIT_33) &
                                                  To_StdLogicVector(INIT_32) &
                                                  To_StdLogicVector(INIT_31) &
                                                  To_StdLogicVector(INIT_30) &
						  To_StdLogicVector(INIT_2F) &
                                                  To_StdLogicVector(INIT_2E) &
                                                  To_StdLogicVector(INIT_2D) &
                                                  To_StdLogicVector(INIT_2C) &
                                                  To_StdLogicVector(INIT_2B) &
                                                  To_StdLogicVector(INIT_2A) &
                                                  To_StdLogicVector(INIT_29) &
                                                  To_StdLogicVector(INIT_28) &
                                                  To_StdLogicVector(INIT_27) &
                                                  To_StdLogicVector(INIT_26) &
                                                  To_StdLogicVector(INIT_25) &
                                                  To_StdLogicVector(INIT_24) &
                                                  To_StdLogicVector(INIT_23) &
                                                  To_StdLogicVector(INIT_22) &
                                                  To_StdLogicVector(INIT_21) &
                                                  To_StdLogicVector(INIT_20) &
						  To_StdLogicVector(INIT_1F) &
                                                  To_StdLogicVector(INIT_1E) &
                                                  To_StdLogicVector(INIT_1D) &
                                                  To_StdLogicVector(INIT_1C) &
                                                  To_StdLogicVector(INIT_1B) &
                                                  To_StdLogicVector(INIT_1A) &
                                                  To_StdLogicVector(INIT_19) &
                                                  To_StdLogicVector(INIT_18) &
                                                  To_StdLogicVector(INIT_17) &
                                                  To_StdLogicVector(INIT_16) &
                                                  To_StdLogicVector(INIT_15) &
                                                  To_StdLogicVector(INIT_14) &
                                                  To_StdLogicVector(INIT_13) &
                                                  To_StdLogicVector(INIT_12) &
                                                  To_StdLogicVector(INIT_11) &
                                                  To_StdLogicVector(INIT_10) & 
						  To_StdLogicVector(INIT_F)  &
                                                  To_StdLogicVector(INIT_E)  &
                                                  To_StdLogicVector(INIT_D)  &
                                                  To_StdLogicVector(INIT_C)  &
                                                  To_StdLogicVector(INIT_B)  &
                                                  To_StdLogicVector(INIT_A)  &
                                                  To_StdLogicVector(INIT_9)  &
                                                  To_StdLogicVector(INIT_8)  &
                                                  To_StdLogicVector(INIT_7)  &
                                                  To_StdLogicVector(INIT_6)  &
                                                  To_StdLogicVector(INIT_5)  &
                                                  To_StdLogicVector(INIT_4)  &
                                                  To_StdLogicVector(INIT_3)  &
                                                  To_StdLogicVector(INIT_2)  &
                                                  To_StdLogicVector(INIT_1)  & 
                                                  To_StdLogicVector(INIT_0) ;  
  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLK'event and (WCLK = '1') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 15 loop
         if (MASK(i) = '0') then
            MEM_temp(16*WADDR_in + i )  := WDATA(i) ;
         end if ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;

  end process ;


  ReadBehavior : process(RCLKN)
  
    variable RADDR_in : integer range 0 to 1023 ;
    variable RDATA_temp : std_logic_vector( 15  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLKN'event and (RCLKN = '0') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 15 loop
            RDATA_temp(i ) := MEM(16*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;

  end process ;

end SB_RAM1024x16NR_ARCH;   --- SB_RAM1024x16NR


---------------------------------------
	--- SB_RAM1024x16NW
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM1024x16NW is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";

           INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";

           INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";

           INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 15  downto 0) ;
                RCLK  : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'H';
                RADDR : in  std_logic_vector( 9  downto 0) ;
                WCLKN : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'H';
                WADDR : in  std_logic_vector( 9  downto 0) ;
                MASK  : in  std_logic_vector( 15  downto 0) ;
                WDATA : in  std_logic_vector( 15  downto 0)
               );
  
  
end SB_RAM1024x16NW;

architecture SB_RAM1024x16NW_ARCH of SB_RAM1024x16NW is

  signal MEM : std_logic_vector(16383 downto 0) ;
  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLKN)
  variable WADDR_in : integer range 0 to 1023;

    variable MEM_temp : std_logic_vector(16383 downto 0) :=  To_StdLogicVector(INIT_3F) &
                                                  To_StdLogicVector(INIT_3E) &
                                                  To_StdLogicVector(INIT_3D) &
                                                  To_StdLogicVector(INIT_3C) &
                                                  To_StdLogicVector(INIT_3B) &
                                                  To_StdLogicVector(INIT_3A) &
                                                  To_StdLogicVector(INIT_39) &
                                                  To_StdLogicVector(INIT_38) &
                                                  To_StdLogicVector(INIT_37) &
                                                  To_StdLogicVector(INIT_36) &
                                                  To_StdLogicVector(INIT_35) &
                                                  To_StdLogicVector(INIT_34) &
                                                  To_StdLogicVector(INIT_33) &
                                                  To_StdLogicVector(INIT_32) &
                                                  To_StdLogicVector(INIT_31) &
                                                  To_StdLogicVector(INIT_30) &
						  To_StdLogicVector(INIT_2F) &
                                                  To_StdLogicVector(INIT_2E) &
                                                  To_StdLogicVector(INIT_2D) &
                                                  To_StdLogicVector(INIT_2C) &
                                                  To_StdLogicVector(INIT_2B) &
                                                  To_StdLogicVector(INIT_2A) &
                                                  To_StdLogicVector(INIT_29) &
                                                  To_StdLogicVector(INIT_28) &
                                                  To_StdLogicVector(INIT_27) &
                                                  To_StdLogicVector(INIT_26) &
                                                  To_StdLogicVector(INIT_25) &
                                                  To_StdLogicVector(INIT_24) &
                                                  To_StdLogicVector(INIT_23) &
                                                  To_StdLogicVector(INIT_22) &
                                                  To_StdLogicVector(INIT_21) &
                                                  To_StdLogicVector(INIT_20) &
						  To_StdLogicVector(INIT_1F) &
                                                  To_StdLogicVector(INIT_1E) &
                                                  To_StdLogicVector(INIT_1D) &
                                                  To_StdLogicVector(INIT_1C) &
                                                  To_StdLogicVector(INIT_1B) &
                                                  To_StdLogicVector(INIT_1A) &
                                                  To_StdLogicVector(INIT_19) &
                                                  To_StdLogicVector(INIT_18) &
                                                  To_StdLogicVector(INIT_17) &
                                                  To_StdLogicVector(INIT_16) &
                                                  To_StdLogicVector(INIT_15) &
                                                  To_StdLogicVector(INIT_14) &
                                                  To_StdLogicVector(INIT_13) &
                                                  To_StdLogicVector(INIT_12) &
                                                  To_StdLogicVector(INIT_11) &
                                                  To_StdLogicVector(INIT_10) & 
						  To_StdLogicVector(INIT_F)  &
                                                  To_StdLogicVector(INIT_E)  &
                                                  To_StdLogicVector(INIT_D)  &
                                                  To_StdLogicVector(INIT_C)  &
                                                  To_StdLogicVector(INIT_B)  &
                                                  To_StdLogicVector(INIT_A)  &
                                                  To_StdLogicVector(INIT_9)  &
                                                  To_StdLogicVector(INIT_8)  &
                                                  To_StdLogicVector(INIT_7)  &
                                                  To_StdLogicVector(INIT_6)  &
                                                  To_StdLogicVector(INIT_5)  &
                                                  To_StdLogicVector(INIT_4)  &
                                                  To_StdLogicVector(INIT_3)  &
                                                  To_StdLogicVector(INIT_2)  &
                                                  To_StdLogicVector(INIT_1)  & 
                                                  To_StdLogicVector(INIT_0) ;  
  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLKN'event and (WCLKN = '0') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 15 loop
         if (MASK(i) = '0') then
            MEM_temp(16*WADDR_in + i )  := WDATA(i) ;
         end if ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;

  end process ;


  ReadBehavior : process(RCLK)
  
    variable RADDR_in : integer range 0 to 1023 ;
    variable RDATA_temp : std_logic_vector( 15  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLK'event and (RCLK = '1') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 15 loop
            RDATA_temp(i ) := MEM(16*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;

  end process ;
 
end SB_RAM1024x16NW_ARCH;   --- SB_RAM1024x16NW



---------------------------------------
	--- SB_RAM1024x16NRNW
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM1024x16NRNW is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";

           INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";

           INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";

           INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 15  downto 0) ;
                RCLKN : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'H';
                RADDR : in  std_logic_vector( 9  downto 0) ;
                WCLKN : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'H';
                WADDR : in  std_logic_vector( 9  downto 0) ;
                MASK  : in  std_logic_vector( 15  downto 0) ;
                WDATA : in  std_logic_vector( 15  downto 0)
               );
  
  
end SB_RAM1024x16NRNW;

architecture SB_RAM1024x16NRNW_ARCH of SB_RAM1024x16NRNW is
 
  signal MEM : std_logic_vector(16383 downto 0) ;
  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLKN)
  variable WADDR_in : integer range 0 to 1023;

    variable MEM_temp : std_logic_vector(16383 downto 0) :=  To_StdLogicVector(INIT_3F) &
                                                  To_StdLogicVector(INIT_3E) &
                                                  To_StdLogicVector(INIT_3D) &
                                                  To_StdLogicVector(INIT_3C) &
                                                  To_StdLogicVector(INIT_3B) &
                                                  To_StdLogicVector(INIT_3A) &
                                                  To_StdLogicVector(INIT_39) &
                                                  To_StdLogicVector(INIT_38) &
                                                  To_StdLogicVector(INIT_37) &
                                                  To_StdLogicVector(INIT_36) &
                                                  To_StdLogicVector(INIT_35) &
                                                  To_StdLogicVector(INIT_34) &
                                                  To_StdLogicVector(INIT_33) &
                                                  To_StdLogicVector(INIT_32) &
                                                  To_StdLogicVector(INIT_31) &
                                                  To_StdLogicVector(INIT_30) &
						  To_StdLogicVector(INIT_2F) &
                                                  To_StdLogicVector(INIT_2E) &
                                                  To_StdLogicVector(INIT_2D) &
                                                  To_StdLogicVector(INIT_2C) &
                                                  To_StdLogicVector(INIT_2B) &
                                                  To_StdLogicVector(INIT_2A) &
                                                  To_StdLogicVector(INIT_29) &
                                                  To_StdLogicVector(INIT_28) &
                                                  To_StdLogicVector(INIT_27) &
                                                  To_StdLogicVector(INIT_26) &
                                                  To_StdLogicVector(INIT_25) &
                                                  To_StdLogicVector(INIT_24) &
                                                  To_StdLogicVector(INIT_23) &
                                                  To_StdLogicVector(INIT_22) &
                                                  To_StdLogicVector(INIT_21) &
                                                  To_StdLogicVector(INIT_20) &
						  To_StdLogicVector(INIT_1F) &
                                                  To_StdLogicVector(INIT_1E) &
                                                  To_StdLogicVector(INIT_1D) &
                                                  To_StdLogicVector(INIT_1C) &
                                                  To_StdLogicVector(INIT_1B) &
                                                  To_StdLogicVector(INIT_1A) &
                                                  To_StdLogicVector(INIT_19) &
                                                  To_StdLogicVector(INIT_18) &
                                                  To_StdLogicVector(INIT_17) &
                                                  To_StdLogicVector(INIT_16) &
                                                  To_StdLogicVector(INIT_15) &
                                                  To_StdLogicVector(INIT_14) &
                                                  To_StdLogicVector(INIT_13) &
                                                  To_StdLogicVector(INIT_12) &
                                                  To_StdLogicVector(INIT_11) &
                                                  To_StdLogicVector(INIT_10) & 
						  To_StdLogicVector(INIT_F)  &
                                                  To_StdLogicVector(INIT_E)  &
                                                  To_StdLogicVector(INIT_D)  &
                                                  To_StdLogicVector(INIT_C)  &
                                                  To_StdLogicVector(INIT_B)  &
                                                  To_StdLogicVector(INIT_A)  &
                                                  To_StdLogicVector(INIT_9)  &
                                                  To_StdLogicVector(INIT_8)  &
                                                  To_StdLogicVector(INIT_7)  &
                                                  To_StdLogicVector(INIT_6)  &
                                                  To_StdLogicVector(INIT_5)  &
                                                  To_StdLogicVector(INIT_4)  &
                                                  To_StdLogicVector(INIT_3)  &
                                                  To_StdLogicVector(INIT_2)  &
                                                  To_StdLogicVector(INIT_1)  & 
                                                  To_StdLogicVector(INIT_0) ;  
  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLKN'event and (WCLKN = '0') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 15 loop
         if (MASK(i) = '0') then
            MEM_temp(16*WADDR_in + i )  := WDATA(i) ;
         end if ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;

  end process ;


  ReadBehavior : process(RCLKN)
  
    variable RADDR_in : integer range 0 to 1023 ;
    variable RDATA_temp : std_logic_vector( 15  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLKN'event and (RCLKN = '0') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 15 loop
            RDATA_temp(i ) := MEM(16*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;
  
end process ;

end SB_RAM1024x16NRNW_ARCH;   --- SB_RAM1024x16NRNW


---------------------------------------
	--- SB_RAM2048x8
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM2048x8 is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";

           INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";

           INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";

           INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 7  downto 0) ;
                RCLK  : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'H';
                RADDR : in  std_logic_vector( 10  downto 0) ;
                WCLK  : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'H';
                WADDR : in  std_logic_vector( 10  downto 0) ;
                WDATA : in  std_logic_vector( 7  downto 0)
               );
  
  
end SB_RAM2048x8;

architecture SB_RAM2048x8_ARCH of SB_RAM2048x8 is

  signal MEM : std_logic_vector(16383 downto 0) ;
  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLK)

    variable WADDR_in : integer range 0 to 2047 ;
    variable MEM_temp : std_logic_vector(16383 downto 0) :=  To_StdLogicVector(INIT_3F) &
                                                  To_StdLogicVector(INIT_3E) &
                                                  To_StdLogicVector(INIT_3D) &
                                                  To_StdLogicVector(INIT_3C) &
                                                  To_StdLogicVector(INIT_3B) &
                                                  To_StdLogicVector(INIT_3A) &
                                                  To_StdLogicVector(INIT_39) &
                                                  To_StdLogicVector(INIT_38) &
                                                  To_StdLogicVector(INIT_37) &
                                                  To_StdLogicVector(INIT_36) &
                                                  To_StdLogicVector(INIT_35) &
                                                  To_StdLogicVector(INIT_34) &
                                                  To_StdLogicVector(INIT_33) &
                                                  To_StdLogicVector(INIT_32) &
                                                  To_StdLogicVector(INIT_31) &
                                                  To_StdLogicVector(INIT_30) &
						  To_StdLogicVector(INIT_2F) &
                                                  To_StdLogicVector(INIT_2E) &
                                                  To_StdLogicVector(INIT_2D) &
                                                  To_StdLogicVector(INIT_2C) &
                                                  To_StdLogicVector(INIT_2B) &
                                                  To_StdLogicVector(INIT_2A) &
                                                  To_StdLogicVector(INIT_29) &
                                                  To_StdLogicVector(INIT_28) &
                                                  To_StdLogicVector(INIT_27) &
                                                  To_StdLogicVector(INIT_26) &
                                                  To_StdLogicVector(INIT_25) &
                                                  To_StdLogicVector(INIT_24) &
                                                  To_StdLogicVector(INIT_23) &
                                                  To_StdLogicVector(INIT_22) &
                                                  To_StdLogicVector(INIT_21) &
                                                  To_StdLogicVector(INIT_20) &
						  To_StdLogicVector(INIT_1F) &
                                                  To_StdLogicVector(INIT_1E) &
                                                  To_StdLogicVector(INIT_1D) &
                                                  To_StdLogicVector(INIT_1C) &
                                                  To_StdLogicVector(INIT_1B) &
                                                  To_StdLogicVector(INIT_1A) &
                                                  To_StdLogicVector(INIT_19) &
                                                  To_StdLogicVector(INIT_18) &
                                                  To_StdLogicVector(INIT_17) &
                                                  To_StdLogicVector(INIT_16) &
                                                  To_StdLogicVector(INIT_15) &
                                                  To_StdLogicVector(INIT_14) &
                                                  To_StdLogicVector(INIT_13) &
                                                  To_StdLogicVector(INIT_12) &
                                                  To_StdLogicVector(INIT_11) &
                                                  To_StdLogicVector(INIT_10) & 
						  To_StdLogicVector(INIT_F)  &
                                                  To_StdLogicVector(INIT_E)  &
                                                  To_StdLogicVector(INIT_D)  &
                                                  To_StdLogicVector(INIT_C)  &
                                                  To_StdLogicVector(INIT_B)  &
                                                  To_StdLogicVector(INIT_A)  &
                                                  To_StdLogicVector(INIT_9)  &
                                                  To_StdLogicVector(INIT_8)  &
                                                  To_StdLogicVector(INIT_7)  &
                                                  To_StdLogicVector(INIT_6)  &
                                                  To_StdLogicVector(INIT_5)  &
                                                  To_StdLogicVector(INIT_4)  &
                                                  To_StdLogicVector(INIT_3)  &
                                                  To_StdLogicVector(INIT_2)  &
                                                  To_StdLogicVector(INIT_1)  & 
                                                  To_StdLogicVector(INIT_0) ;  

  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLK'event and (WCLK = '1') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 7 loop
            MEM_temp(8*WADDR_in + i )  := WDATA(i) ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;


  end process ;


  ReadBehavior : process(RCLK)
  
    variable RADDR_in : integer range 0 to 2047 ;
    variable RDATA_temp : std_logic_vector( 7  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLK'event and (RCLK = '1') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 7 loop
            RDATA_temp(i ) := MEM(8*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;

  end process ;

end SB_RAM2048x8_ARCH;   --- SB_RAM2048x8

---------------------------------------
	--- SB_RAM2048x8NR
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM2048x8NR is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";

           INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";

           INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";

           INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 7  downto 0) ;
                RCLKN : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'H';
                RADDR : in  std_logic_vector( 10  downto 0) ;
                WCLK  : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'H';
                WADDR : in  std_logic_vector( 10  downto 0) ;
                WDATA : in  std_logic_vector( 7  downto 0)
               );
  
  
end SB_RAM2048x8NR;

architecture SB_RAM2048x8NR_ARCH of SB_RAM2048x8NR is

  signal MEM : std_logic_vector(16383 downto 0) ;
  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLK)

    variable WADDR_in : integer range 0 to 2047 ;
    variable MEM_temp : std_logic_vector(16383 downto 0) :=  To_StdLogicVector(INIT_3F) &
                                                  To_StdLogicVector(INIT_3E) &
                                                  To_StdLogicVector(INIT_3D) &
                                                  To_StdLogicVector(INIT_3C) &
                                                  To_StdLogicVector(INIT_3B) &
                                                  To_StdLogicVector(INIT_3A) &
                                                  To_StdLogicVector(INIT_39) &
                                                  To_StdLogicVector(INIT_38) &
                                                  To_StdLogicVector(INIT_37) &
                                                  To_StdLogicVector(INIT_36) &
                                                  To_StdLogicVector(INIT_35) &
                                                  To_StdLogicVector(INIT_34) &
                                                  To_StdLogicVector(INIT_33) &
                                                  To_StdLogicVector(INIT_32) &
                                                  To_StdLogicVector(INIT_31) &
                                                  To_StdLogicVector(INIT_30) &
						  To_StdLogicVector(INIT_2F) &
                                                  To_StdLogicVector(INIT_2E) &
                                                  To_StdLogicVector(INIT_2D) &
                                                  To_StdLogicVector(INIT_2C) &
                                                  To_StdLogicVector(INIT_2B) &
                                                  To_StdLogicVector(INIT_2A) &
                                                  To_StdLogicVector(INIT_29) &
                                                  To_StdLogicVector(INIT_28) &
                                                  To_StdLogicVector(INIT_27) &
                                                  To_StdLogicVector(INIT_26) &
                                                  To_StdLogicVector(INIT_25) &
                                                  To_StdLogicVector(INIT_24) &
                                                  To_StdLogicVector(INIT_23) &
                                                  To_StdLogicVector(INIT_22) &
                                                  To_StdLogicVector(INIT_21) &
                                                  To_StdLogicVector(INIT_20) &
						  To_StdLogicVector(INIT_1F) &
                                                  To_StdLogicVector(INIT_1E) &
                                                  To_StdLogicVector(INIT_1D) &
                                                  To_StdLogicVector(INIT_1C) &
                                                  To_StdLogicVector(INIT_1B) &
                                                  To_StdLogicVector(INIT_1A) &
                                                  To_StdLogicVector(INIT_19) &
                                                  To_StdLogicVector(INIT_18) &
                                                  To_StdLogicVector(INIT_17) &
                                                  To_StdLogicVector(INIT_16) &
                                                  To_StdLogicVector(INIT_15) &
                                                  To_StdLogicVector(INIT_14) &
                                                  To_StdLogicVector(INIT_13) &
                                                  To_StdLogicVector(INIT_12) &
                                                  To_StdLogicVector(INIT_11) &
                                                  To_StdLogicVector(INIT_10) & 
						  To_StdLogicVector(INIT_F)  &
                                                  To_StdLogicVector(INIT_E)  &
                                                  To_StdLogicVector(INIT_D)  &
                                                  To_StdLogicVector(INIT_C)  &
                                                  To_StdLogicVector(INIT_B)  &
                                                  To_StdLogicVector(INIT_A)  &
                                                  To_StdLogicVector(INIT_9)  &
                                                  To_StdLogicVector(INIT_8)  &
                                                  To_StdLogicVector(INIT_7)  &
                                                  To_StdLogicVector(INIT_6)  &
                                                  To_StdLogicVector(INIT_5)  &
                                                  To_StdLogicVector(INIT_4)  &
                                                  To_StdLogicVector(INIT_3)  &
                                                  To_StdLogicVector(INIT_2)  &
                                                  To_StdLogicVector(INIT_1)  & 
                                                  To_StdLogicVector(INIT_0) ;  

  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLK'event and (WCLK = '1') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 7 loop
            MEM_temp(8*WADDR_in + i )  := WDATA(i) ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;


  end process ;


  ReadBehavior : process(RCLKN)
  
    variable RADDR_in : integer range 0 to 2047 ;
    variable RDATA_temp : std_logic_vector( 7  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLKN'event and (RCLKN = '0') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 7 loop
            RDATA_temp(i ) := MEM(8*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;

  end process ;

end SB_RAM2048x8NR_ARCH;   --- SB_RAM2048x8NR



---------------------------------------
	--- SB_RAM2048x8NW
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM2048x8NW is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";

           INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";

           INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 7  downto 0) ;
                RCLK  : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'H';
                RADDR : in  std_logic_vector( 10  downto 0) ;
                WCLKN : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'H';
                WADDR : in  std_logic_vector( 10  downto 0) ;
                WDATA : in  std_logic_vector( 7  downto 0)
               );
  
  
end SB_RAM2048x8NW;

architecture SB_RAM2048x8NW_ARCH of SB_RAM2048x8NW is

  signal MEM : std_logic_vector(16383 downto 0) ;
  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLKN)

    variable WADDR_in : integer range 0 to 2047 ;
    variable MEM_temp : std_logic_vector(16383 downto 0) :=  To_StdLogicVector(INIT_3F) &
                                                  To_StdLogicVector(INIT_3E) &
                                                  To_StdLogicVector(INIT_3D) &
                                                  To_StdLogicVector(INIT_3C) &
                                                  To_StdLogicVector(INIT_3B) &
                                                  To_StdLogicVector(INIT_3A) &
                                                  To_StdLogicVector(INIT_39) &
                                                  To_StdLogicVector(INIT_38) &
                                                  To_StdLogicVector(INIT_37) &
                                                  To_StdLogicVector(INIT_36) &
                                                  To_StdLogicVector(INIT_35) &
                                                  To_StdLogicVector(INIT_34) &
                                                  To_StdLogicVector(INIT_33) &
                                                  To_StdLogicVector(INIT_32) &
                                                  To_StdLogicVector(INIT_31) &
                                                  To_StdLogicVector(INIT_30) &
						  To_StdLogicVector(INIT_2F) &
                                                  To_StdLogicVector(INIT_2E) &
                                                  To_StdLogicVector(INIT_2D) &
                                                  To_StdLogicVector(INIT_2C) &
                                                  To_StdLogicVector(INIT_2B) &
                                                  To_StdLogicVector(INIT_2A) &
                                                  To_StdLogicVector(INIT_29) &
                                                  To_StdLogicVector(INIT_28) &
                                                  To_StdLogicVector(INIT_27) &
                                                  To_StdLogicVector(INIT_26) &
                                                  To_StdLogicVector(INIT_25) &
                                                  To_StdLogicVector(INIT_24) &
                                                  To_StdLogicVector(INIT_23) &
                                                  To_StdLogicVector(INIT_22) &
                                                  To_StdLogicVector(INIT_21) &
                                                  To_StdLogicVector(INIT_20) &
						  To_StdLogicVector(INIT_1F) &
                                                  To_StdLogicVector(INIT_1E) &
                                                  To_StdLogicVector(INIT_1D) &
                                                  To_StdLogicVector(INIT_1C) &
                                                  To_StdLogicVector(INIT_1B) &
                                                  To_StdLogicVector(INIT_1A) &
                                                  To_StdLogicVector(INIT_19) &
                                                  To_StdLogicVector(INIT_18) &
                                                  To_StdLogicVector(INIT_17) &
                                                  To_StdLogicVector(INIT_16) &
                                                  To_StdLogicVector(INIT_15) &
                                                  To_StdLogicVector(INIT_14) &
                                                  To_StdLogicVector(INIT_13) &
                                                  To_StdLogicVector(INIT_12) &
                                                  To_StdLogicVector(INIT_11) &
                                                  To_StdLogicVector(INIT_10) & 
						  To_StdLogicVector(INIT_F)  &
                                                  To_StdLogicVector(INIT_E)  &
                                                  To_StdLogicVector(INIT_D)  &
                                                  To_StdLogicVector(INIT_C)  &
                                                  To_StdLogicVector(INIT_B)  &
                                                  To_StdLogicVector(INIT_A)  &
                                                  To_StdLogicVector(INIT_9)  &
                                                  To_StdLogicVector(INIT_8)  &
                                                  To_StdLogicVector(INIT_7)  &
                                                  To_StdLogicVector(INIT_6)  &
                                                  To_StdLogicVector(INIT_5)  &
                                                  To_StdLogicVector(INIT_4)  &
                                                  To_StdLogicVector(INIT_3)  &
                                                  To_StdLogicVector(INIT_2)  &
                                                  To_StdLogicVector(INIT_1)  & 
                                                  To_StdLogicVector(INIT_0) ;  

  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLKN'event and (WCLKN = '0') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 7 loop
            MEM_temp(8*WADDR_in + i )  := WDATA(i) ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;


  end process ;


  ReadBehavior : process(RCLK)
  
    variable RADDR_in : integer range 0 to 2047 ;
    variable RDATA_temp : std_logic_vector( 7  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLK'event and (RCLK = '1') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 7 loop
            RDATA_temp(i ) := MEM(8*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;

  end process ;

end SB_RAM2048x8NW_ARCH;   --- SB_RAM2048x8NW


---------------------------------------
	--- SB_RAM2048x8NRNW
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM2048x8NRNW is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 7  downto 0) ;
                RCLKN : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'H';
                RADDR : in  std_logic_vector( 10  downto 0) ;
                WCLKN : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'H';
                WADDR : in  std_logic_vector( 10  downto 0) ;
                WDATA : in  std_logic_vector( 7  downto 0)
               );
  
  
end SB_RAM2048x8NRNW;

architecture SB_RAM2048x8NRNW_ARCH of SB_RAM2048x8NRNW is
 
  signal MEM : std_logic_vector(16383 downto 0) ;
  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLKN)

    variable WADDR_in : integer range 0 to 2047 ;
    variable MEM_temp : std_logic_vector(16383 downto 0) :=  To_StdLogicVector(INIT_3F) &
                                                  To_StdLogicVector(INIT_3E) &
                                                  To_StdLogicVector(INIT_3D) &
                                                  To_StdLogicVector(INIT_3C) &
                                                  To_StdLogicVector(INIT_3B) &
                                                  To_StdLogicVector(INIT_3A) &
                                                  To_StdLogicVector(INIT_39) &
                                                  To_StdLogicVector(INIT_38) &
                                                  To_StdLogicVector(INIT_37) &
                                                  To_StdLogicVector(INIT_36) &
                                                  To_StdLogicVector(INIT_35) &
                                                  To_StdLogicVector(INIT_34) &
                                                  To_StdLogicVector(INIT_33) &
                                                  To_StdLogicVector(INIT_32) &
                                                  To_StdLogicVector(INIT_31) &
                                                  To_StdLogicVector(INIT_30) &
						  To_StdLogicVector(INIT_2F) &
                                                  To_StdLogicVector(INIT_2E) &
                                                  To_StdLogicVector(INIT_2D) &
                                                  To_StdLogicVector(INIT_2C) &
                                                  To_StdLogicVector(INIT_2B) &
                                                  To_StdLogicVector(INIT_2A) &
                                                  To_StdLogicVector(INIT_29) &
                                                  To_StdLogicVector(INIT_28) &
                                                  To_StdLogicVector(INIT_27) &
                                                  To_StdLogicVector(INIT_26) &
                                                  To_StdLogicVector(INIT_25) &
                                                  To_StdLogicVector(INIT_24) &
                                                  To_StdLogicVector(INIT_23) &
                                                  To_StdLogicVector(INIT_22) &
                                                  To_StdLogicVector(INIT_21) &
                                                  To_StdLogicVector(INIT_20) &
						  To_StdLogicVector(INIT_1F) &
                                                  To_StdLogicVector(INIT_1E) &
                                                  To_StdLogicVector(INIT_1D) &
                                                  To_StdLogicVector(INIT_1C) &
                                                  To_StdLogicVector(INIT_1B) &
                                                  To_StdLogicVector(INIT_1A) &
                                                  To_StdLogicVector(INIT_19) &
                                                  To_StdLogicVector(INIT_18) &
                                                  To_StdLogicVector(INIT_17) &
                                                  To_StdLogicVector(INIT_16) &
                                                  To_StdLogicVector(INIT_15) &
                                                  To_StdLogicVector(INIT_14) &
                                                  To_StdLogicVector(INIT_13) &
                                                  To_StdLogicVector(INIT_12) &
                                                  To_StdLogicVector(INIT_11) &
                                                  To_StdLogicVector(INIT_10) & 
						  To_StdLogicVector(INIT_F)  &
                                                  To_StdLogicVector(INIT_E)  &
                                                  To_StdLogicVector(INIT_D)  &
                                                  To_StdLogicVector(INIT_C)  &
                                                  To_StdLogicVector(INIT_B)  &
                                                  To_StdLogicVector(INIT_A)  &
                                                  To_StdLogicVector(INIT_9)  &
                                                  To_StdLogicVector(INIT_8)  &
                                                  To_StdLogicVector(INIT_7)  &
                                                  To_StdLogicVector(INIT_6)  &
                                                  To_StdLogicVector(INIT_5)  &
                                                  To_StdLogicVector(INIT_4)  &
                                                  To_StdLogicVector(INIT_3)  &
                                                  To_StdLogicVector(INIT_2)  &
                                                  To_StdLogicVector(INIT_1)  & 
                                                  To_StdLogicVector(INIT_0) ;  

  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLKN'event and (WCLKN = '0') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 7 loop
            MEM_temp(8*WADDR_in + i )  := WDATA(i) ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;


  end process ;


  ReadBehavior : process(RCLKN)
  
    variable RADDR_in : integer range 0 to 2047 ;
    variable RDATA_temp : std_logic_vector( 7  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLKN'event and (RCLKN = '0') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 7 loop
            RDATA_temp(i ) := MEM(8*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;

  end process ;

end SB_RAM2048x8NRNW_ARCH;   --- SB_RAM2048x8NRNW


---------------------------------------
	--- SB_RAM4096x4
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM4096x4 is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 3  downto 0) ;
                RCLK  : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'H';
                RADDR : in  std_logic_vector( 11  downto 0) ;
                WCLK  : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'H';
                WADDR : in  std_logic_vector( 11  downto 0) ;
                WDATA : in  std_logic_vector( 3  downto 0)
               );
  
  
end SB_RAM4096x4;

architecture SB_RAM4096x4_ARCH of SB_RAM4096x4 is

  signal MEM : std_logic_vector(16383 downto 0) ;
  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLK)
    variable WADDR_in : integer range 0 to 4095 ;
    variable MEM_temp : std_logic_vector(16383 downto 0) :=  To_StdLogicVector(INIT_3F) &
                                                  To_StdLogicVector(INIT_3E) &
                                                  To_StdLogicVector(INIT_3D) &
                                                  To_StdLogicVector(INIT_3C) &
                                                  To_StdLogicVector(INIT_3B) &
                                                  To_StdLogicVector(INIT_3A) &
                                                  To_StdLogicVector(INIT_39) &
                                                  To_StdLogicVector(INIT_38) &
                                                  To_StdLogicVector(INIT_37) &
                                                  To_StdLogicVector(INIT_36) &
                                                  To_StdLogicVector(INIT_35) &
                                                  To_StdLogicVector(INIT_34) &
                                                  To_StdLogicVector(INIT_33) &
                                                  To_StdLogicVector(INIT_32) &
                                                  To_StdLogicVector(INIT_31) &
                                                  To_StdLogicVector(INIT_30) &
						  To_StdLogicVector(INIT_2F) &
                                                  To_StdLogicVector(INIT_2E) &
                                                  To_StdLogicVector(INIT_2D) &
                                                  To_StdLogicVector(INIT_2C) &
                                                  To_StdLogicVector(INIT_2B) &
                                                  To_StdLogicVector(INIT_2A) &
                                                  To_StdLogicVector(INIT_29) &
                                                  To_StdLogicVector(INIT_28) &
                                                  To_StdLogicVector(INIT_27) &
                                                  To_StdLogicVector(INIT_26) &
                                                  To_StdLogicVector(INIT_25) &
                                                  To_StdLogicVector(INIT_24) &
                                                  To_StdLogicVector(INIT_23) &
                                                  To_StdLogicVector(INIT_22) &
                                                  To_StdLogicVector(INIT_21) &
                                                  To_StdLogicVector(INIT_20) &
						  To_StdLogicVector(INIT_1F) &
                                                  To_StdLogicVector(INIT_1E) &
                                                  To_StdLogicVector(INIT_1D) &
                                                  To_StdLogicVector(INIT_1C) &
                                                  To_StdLogicVector(INIT_1B) &
                                                  To_StdLogicVector(INIT_1A) &
                                                  To_StdLogicVector(INIT_19) &
                                                  To_StdLogicVector(INIT_18) &
                                                  To_StdLogicVector(INIT_17) &
                                                  To_StdLogicVector(INIT_16) &
                                                  To_StdLogicVector(INIT_15) &
                                                  To_StdLogicVector(INIT_14) &
                                                  To_StdLogicVector(INIT_13) &
                                                  To_StdLogicVector(INIT_12) &
                                                  To_StdLogicVector(INIT_11) &
                                                  To_StdLogicVector(INIT_10) & 
						  To_StdLogicVector(INIT_F)  &
                                                  To_StdLogicVector(INIT_E)  &
                                                  To_StdLogicVector(INIT_D)  &
                                                  To_StdLogicVector(INIT_C)  &
                                                  To_StdLogicVector(INIT_B)  &
                                                  To_StdLogicVector(INIT_A)  &
                                                  To_StdLogicVector(INIT_9)  &
                                                  To_StdLogicVector(INIT_8)  &
                                                  To_StdLogicVector(INIT_7)  &
                                                  To_StdLogicVector(INIT_6)  &
                                                  To_StdLogicVector(INIT_5)  &
                                                  To_StdLogicVector(INIT_4)  &
                                                  To_StdLogicVector(INIT_3)  &
                                                  To_StdLogicVector(INIT_2)  &
                                                  To_StdLogicVector(INIT_1)  & 
                                                  To_StdLogicVector(INIT_0) ;  

  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLK'event and (WCLK = '1') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 3 loop
            MEM_temp(4*WADDR_in + i )  := WDATA(i) ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;


  end process ;


  ReadBehavior : process(RCLK)
  
    variable RADDR_in : integer range 0 to 4095;
    variable RDATA_temp : std_logic_vector( 3  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLK'event and (RCLK = '1') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 3 loop
            RDATA_temp(i ) := MEM(4*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;

  end process ;

end SB_RAM4096x4_ARCH;   --- SB_RAM4096x4

---------------------------------------
	--- SB_RAM4096x4NR
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM4096x4NR is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 3  downto 0) ;
                RCLKN : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'H';
                RADDR : in  std_logic_vector( 11  downto 0) ;
                WCLK  : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'H';
                WADDR : in  std_logic_vector( 11  downto 0) ;
                WDATA : in  std_logic_vector( 3  downto 0)
               );
  
end SB_RAM4096x4NR;

architecture SB_RAM4096x4NR_ARCH of SB_RAM4096x4NR is

  signal MEM : std_logic_vector(16383 downto 0) ;
  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLK)
    variable WADDR_in : integer range 0 to 4095 ;
    variable MEM_temp : std_logic_vector(16383 downto 0) :=  To_StdLogicVector(INIT_3F) &
                                                  To_StdLogicVector(INIT_3E) &
                                                  To_StdLogicVector(INIT_3D) &
                                                  To_StdLogicVector(INIT_3C) &
                                                  To_StdLogicVector(INIT_3B) &
                                                  To_StdLogicVector(INIT_3A) &
                                                  To_StdLogicVector(INIT_39) &
                                                  To_StdLogicVector(INIT_38) &
                                                  To_StdLogicVector(INIT_37) &
                                                  To_StdLogicVector(INIT_36) &
                                                  To_StdLogicVector(INIT_35) &
                                                  To_StdLogicVector(INIT_34) &
                                                  To_StdLogicVector(INIT_33) &
                                                  To_StdLogicVector(INIT_32) &
                                                  To_StdLogicVector(INIT_31) &
                                                  To_StdLogicVector(INIT_30) &
						  To_StdLogicVector(INIT_2F) &
                                                  To_StdLogicVector(INIT_2E) &
                                                  To_StdLogicVector(INIT_2D) &
                                                  To_StdLogicVector(INIT_2C) &
                                                  To_StdLogicVector(INIT_2B) &
                                                  To_StdLogicVector(INIT_2A) &
                                                  To_StdLogicVector(INIT_29) &
                                                  To_StdLogicVector(INIT_28) &
                                                  To_StdLogicVector(INIT_27) &
                                                  To_StdLogicVector(INIT_26) &
                                                  To_StdLogicVector(INIT_25) &
                                                  To_StdLogicVector(INIT_24) &
                                                  To_StdLogicVector(INIT_23) &
                                                  To_StdLogicVector(INIT_22) &
                                                  To_StdLogicVector(INIT_21) &
                                                  To_StdLogicVector(INIT_20) &
						  To_StdLogicVector(INIT_1F) &
                                                  To_StdLogicVector(INIT_1E) &
                                                  To_StdLogicVector(INIT_1D) &
                                                  To_StdLogicVector(INIT_1C) &
                                                  To_StdLogicVector(INIT_1B) &
                                                  To_StdLogicVector(INIT_1A) &
                                                  To_StdLogicVector(INIT_19) &
                                                  To_StdLogicVector(INIT_18) &
                                                  To_StdLogicVector(INIT_17) &
                                                  To_StdLogicVector(INIT_16) &
                                                  To_StdLogicVector(INIT_15) &
                                                  To_StdLogicVector(INIT_14) &
                                                  To_StdLogicVector(INIT_13) &
                                                  To_StdLogicVector(INIT_12) &
                                                  To_StdLogicVector(INIT_11) &
                                                  To_StdLogicVector(INIT_10) & 
						  To_StdLogicVector(INIT_F)  &
                                                  To_StdLogicVector(INIT_E)  &
                                                  To_StdLogicVector(INIT_D)  &
                                                  To_StdLogicVector(INIT_C)  &
                                                  To_StdLogicVector(INIT_B)  &
                                                  To_StdLogicVector(INIT_A)  &
                                                  To_StdLogicVector(INIT_9)  &
                                                  To_StdLogicVector(INIT_8)  &
                                                  To_StdLogicVector(INIT_7)  &
                                                  To_StdLogicVector(INIT_6)  &
                                                  To_StdLogicVector(INIT_5)  &
                                                  To_StdLogicVector(INIT_4)  &
                                                  To_StdLogicVector(INIT_3)  &
                                                  To_StdLogicVector(INIT_2)  &
                                                  To_StdLogicVector(INIT_1)  & 
                                                  To_StdLogicVector(INIT_0) ;  

  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLK'event and (WCLK = '1') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 3 loop
            MEM_temp(4*WADDR_in + i )  := WDATA(i) ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;


  end process ;


  ReadBehavior : process(RCLKN)
  
    variable RADDR_in : integer range 0 to 4095;
    variable RDATA_temp : std_logic_vector( 3  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLKN'event and (RCLKN = '0') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 3 loop
            RDATA_temp(i ) := MEM(4*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;

  end process ;

end SB_RAM4096x4NR_ARCH;   --- SB_RAM4096x4NR

---------------------------------------
	--- SB_RAM4096x4NW
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM4096x4NW is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 3  downto 0) ;
                RCLK  : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'H';
                RADDR : in  std_logic_vector( 11  downto 0) ;
                WCLKN : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'H';
                WADDR : in  std_logic_vector( 11  downto 0) ;
                WDATA : in  std_logic_vector( 3  downto 0)
               );
  
end SB_RAM4096x4NW;

architecture SB_RAM4096x4NW_ARCH of SB_RAM4096x4NW is
 
  signal MEM : std_logic_vector(16383 downto 0) ;
  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLKN)
    variable WADDR_in : integer range 0 to 4095 ;
    variable MEM_temp : std_logic_vector(16383 downto 0) :=  To_StdLogicVector(INIT_3F) &
                                                  To_StdLogicVector(INIT_3E) &
                                                  To_StdLogicVector(INIT_3D) &
                                                  To_StdLogicVector(INIT_3C) &
                                                  To_StdLogicVector(INIT_3B) &
                                                  To_StdLogicVector(INIT_3A) &
                                                  To_StdLogicVector(INIT_39) &
                                                  To_StdLogicVector(INIT_38) &
                                                  To_StdLogicVector(INIT_37) &
                                                  To_StdLogicVector(INIT_36) &
                                                  To_StdLogicVector(INIT_35) &
                                                  To_StdLogicVector(INIT_34) &
                                                  To_StdLogicVector(INIT_33) &
                                                  To_StdLogicVector(INIT_32) &
                                                  To_StdLogicVector(INIT_31) &
                                                  To_StdLogicVector(INIT_30) &
						  To_StdLogicVector(INIT_2F) &
                                                  To_StdLogicVector(INIT_2E) &
                                                  To_StdLogicVector(INIT_2D) &
                                                  To_StdLogicVector(INIT_2C) &
                                                  To_StdLogicVector(INIT_2B) &
                                                  To_StdLogicVector(INIT_2A) &
                                                  To_StdLogicVector(INIT_29) &
                                                  To_StdLogicVector(INIT_28) &
                                                  To_StdLogicVector(INIT_27) &
                                                  To_StdLogicVector(INIT_26) &
                                                  To_StdLogicVector(INIT_25) &
                                                  To_StdLogicVector(INIT_24) &
                                                  To_StdLogicVector(INIT_23) &
                                                  To_StdLogicVector(INIT_22) &
                                                  To_StdLogicVector(INIT_21) &
                                                  To_StdLogicVector(INIT_20) &
						  To_StdLogicVector(INIT_1F) &
                                                  To_StdLogicVector(INIT_1E) &
                                                  To_StdLogicVector(INIT_1D) &
                                                  To_StdLogicVector(INIT_1C) &
                                                  To_StdLogicVector(INIT_1B) &
                                                  To_StdLogicVector(INIT_1A) &
                                                  To_StdLogicVector(INIT_19) &
                                                  To_StdLogicVector(INIT_18) &
                                                  To_StdLogicVector(INIT_17) &
                                                  To_StdLogicVector(INIT_16) &
                                                  To_StdLogicVector(INIT_15) &
                                                  To_StdLogicVector(INIT_14) &
                                                  To_StdLogicVector(INIT_13) &
                                                  To_StdLogicVector(INIT_12) &
                                                  To_StdLogicVector(INIT_11) &
                                                  To_StdLogicVector(INIT_10) & 
						  To_StdLogicVector(INIT_F)  &
                                                  To_StdLogicVector(INIT_E)  &
                                                  To_StdLogicVector(INIT_D)  &
                                                  To_StdLogicVector(INIT_C)  &
                                                  To_StdLogicVector(INIT_B)  &
                                                  To_StdLogicVector(INIT_A)  &
                                                  To_StdLogicVector(INIT_9)  &
                                                  To_StdLogicVector(INIT_8)  &
                                                  To_StdLogicVector(INIT_7)  &
                                                  To_StdLogicVector(INIT_6)  &
                                                  To_StdLogicVector(INIT_5)  &
                                                  To_StdLogicVector(INIT_4)  &
                                                  To_StdLogicVector(INIT_3)  &
                                                  To_StdLogicVector(INIT_2)  &
                                                  To_StdLogicVector(INIT_1)  & 
                                                  To_StdLogicVector(INIT_0) ;  

  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLKN'event and (WCLKN = '0') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 3 loop
            MEM_temp(4*WADDR_in + i )  := WDATA(i) ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;

  end process ;


  ReadBehavior : process(RCLK)
  
    variable RADDR_in : integer range 0 to 4095;
    variable RDATA_temp : std_logic_vector( 3  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLK'event and (RCLK = '1') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 3 loop
            RDATA_temp(i ) := MEM(4*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;

  end process ;

end SB_RAM4096x4NW_ARCH;   --- SB_RAM4096x4NW


---------------------------------------
	--- SB_RAM4096x4NRNW
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM4096x4NRNW is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 3  downto 0) ;
                RCLKN : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'H';
                RADDR : in  std_logic_vector( 11  downto 0) ;
                WCLKN : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'H';
                WADDR : in  std_logic_vector( 11  downto 0) ;
                WDATA : in  std_logic_vector( 3  downto 0)
               );
  
  
end SB_RAM4096x4NRNW;

architecture SB_RAM4096x4NRNW_ARCH of SB_RAM4096x4NRNW is
 
  signal MEM : std_logic_vector(16383 downto 0) ;
  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLKN)
    variable WADDR_in : integer range 0 to 4095 ;
    variable MEM_temp : std_logic_vector(16383 downto 0) :=  To_StdLogicVector(INIT_3F) &
                                                  To_StdLogicVector(INIT_3E) &
                                                  To_StdLogicVector(INIT_3D) &
                                                  To_StdLogicVector(INIT_3C) &
                                                  To_StdLogicVector(INIT_3B) &
                                                  To_StdLogicVector(INIT_3A) &
                                                  To_StdLogicVector(INIT_39) &
                                                  To_StdLogicVector(INIT_38) &
                                                  To_StdLogicVector(INIT_37) &
                                                  To_StdLogicVector(INIT_36) &
                                                  To_StdLogicVector(INIT_35) &
                                                  To_StdLogicVector(INIT_34) &
                                                  To_StdLogicVector(INIT_33) &
                                                  To_StdLogicVector(INIT_32) &
                                                  To_StdLogicVector(INIT_31) &
                                                  To_StdLogicVector(INIT_30) &
						  To_StdLogicVector(INIT_2F) &
                                                  To_StdLogicVector(INIT_2E) &
                                                  To_StdLogicVector(INIT_2D) &
                                                  To_StdLogicVector(INIT_2C) &
                                                  To_StdLogicVector(INIT_2B) &
                                                  To_StdLogicVector(INIT_2A) &
                                                  To_StdLogicVector(INIT_29) &
                                                  To_StdLogicVector(INIT_28) &
                                                  To_StdLogicVector(INIT_27) &
                                                  To_StdLogicVector(INIT_26) &
                                                  To_StdLogicVector(INIT_25) &
                                                  To_StdLogicVector(INIT_24) &
                                                  To_StdLogicVector(INIT_23) &
                                                  To_StdLogicVector(INIT_22) &
                                                  To_StdLogicVector(INIT_21) &
                                                  To_StdLogicVector(INIT_20) &
						  To_StdLogicVector(INIT_1F) &
                                                  To_StdLogicVector(INIT_1E) &
                                                  To_StdLogicVector(INIT_1D) &
                                                  To_StdLogicVector(INIT_1C) &
                                                  To_StdLogicVector(INIT_1B) &
                                                  To_StdLogicVector(INIT_1A) &
                                                  To_StdLogicVector(INIT_19) &
                                                  To_StdLogicVector(INIT_18) &
                                                  To_StdLogicVector(INIT_17) &
                                                  To_StdLogicVector(INIT_16) &
                                                  To_StdLogicVector(INIT_15) &
                                                  To_StdLogicVector(INIT_14) &
                                                  To_StdLogicVector(INIT_13) &
                                                  To_StdLogicVector(INIT_12) &
                                                  To_StdLogicVector(INIT_11) &
                                                  To_StdLogicVector(INIT_10) & 
						  To_StdLogicVector(INIT_F)  &
                                                  To_StdLogicVector(INIT_E)  &
                                                  To_StdLogicVector(INIT_D)  &
                                                  To_StdLogicVector(INIT_C)  &
                                                  To_StdLogicVector(INIT_B)  &
                                                  To_StdLogicVector(INIT_A)  &
                                                  To_StdLogicVector(INIT_9)  &
                                                  To_StdLogicVector(INIT_8)  &
                                                  To_StdLogicVector(INIT_7)  &
                                                  To_StdLogicVector(INIT_6)  &
                                                  To_StdLogicVector(INIT_5)  &
                                                  To_StdLogicVector(INIT_4)  &
                                                  To_StdLogicVector(INIT_3)  &
                                                  To_StdLogicVector(INIT_2)  &
                                                  To_StdLogicVector(INIT_1)  & 
                                                  To_StdLogicVector(INIT_0) ;  

  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLKN'event and (WCLKN = '0') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 3 loop
            MEM_temp(4*WADDR_in + i )  := WDATA(i) ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;


  end process ;


  ReadBehavior : process(RCLKN)
  
    variable RADDR_in : integer range 0 to 4095;
    variable RDATA_temp : std_logic_vector( 3  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLKN'event and (RCLKN = '0') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 3 loop
            RDATA_temp(i ) := MEM(4*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;

  end process ;

end SB_RAM4096x4NRNW_ARCH;   --- SB_RAM4096x4NRNW


---------------------------------------
	--- SB_RAM8192x2
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM8192x2 is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 1  downto 0) ;
                RCLK  : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'H';
                RADDR : in  std_logic_vector( 12  downto 0) ;
                WCLK  : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'H';
                WADDR : in  std_logic_vector( 12  downto 0) ;
                WDATA : in  std_logic_vector( 1  downto 0)
               );
  
  
end SB_RAM8192x2;

architecture SB_RAM8192x2_ARCH of SB_RAM8192x2 is

  signal MEM : std_logic_vector(16383 downto 0) ;
  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLK)
    variable WADDR_in : integer range 0 to 8191;
    variable MEM_temp : std_logic_vector(16383 downto 0) :=  To_StdLogicVector(INIT_3F) &
                                                  To_StdLogicVector(INIT_3E) &
                                                  To_StdLogicVector(INIT_3D) &
                                                  To_StdLogicVector(INIT_3C) &
                                                  To_StdLogicVector(INIT_3B) &
                                                  To_StdLogicVector(INIT_3A) &
                                                  To_StdLogicVector(INIT_39) &
                                                  To_StdLogicVector(INIT_38) &
                                                  To_StdLogicVector(INIT_37) &
                                                  To_StdLogicVector(INIT_36) &
                                                  To_StdLogicVector(INIT_35) &
                                                  To_StdLogicVector(INIT_34) &
                                                  To_StdLogicVector(INIT_33) &
                                                  To_StdLogicVector(INIT_32) &
                                                  To_StdLogicVector(INIT_31) &
                                                  To_StdLogicVector(INIT_30) &
						  To_StdLogicVector(INIT_2F) &
                                                  To_StdLogicVector(INIT_2E) &
                                                  To_StdLogicVector(INIT_2D) &
                                                  To_StdLogicVector(INIT_2C) &
                                                  To_StdLogicVector(INIT_2B) &
                                                  To_StdLogicVector(INIT_2A) &
                                                  To_StdLogicVector(INIT_29) &
                                                  To_StdLogicVector(INIT_28) &
                                                  To_StdLogicVector(INIT_27) &
                                                  To_StdLogicVector(INIT_26) &
                                                  To_StdLogicVector(INIT_25) &
                                                  To_StdLogicVector(INIT_24) &
                                                  To_StdLogicVector(INIT_23) &
                                                  To_StdLogicVector(INIT_22) &
                                                  To_StdLogicVector(INIT_21) &
                                                  To_StdLogicVector(INIT_20) &
						  To_StdLogicVector(INIT_1F) &
                                                  To_StdLogicVector(INIT_1E) &
                                                  To_StdLogicVector(INIT_1D) &
                                                  To_StdLogicVector(INIT_1C) &
                                                  To_StdLogicVector(INIT_1B) &
                                                  To_StdLogicVector(INIT_1A) &
                                                  To_StdLogicVector(INIT_19) &
                                                  To_StdLogicVector(INIT_18) &
                                                  To_StdLogicVector(INIT_17) &
                                                  To_StdLogicVector(INIT_16) &
                                                  To_StdLogicVector(INIT_15) &
                                                  To_StdLogicVector(INIT_14) &
                                                  To_StdLogicVector(INIT_13) &
                                                  To_StdLogicVector(INIT_12) &
                                                  To_StdLogicVector(INIT_11) &
                                                  To_StdLogicVector(INIT_10) & 
						  To_StdLogicVector(INIT_F)  &
                                                  To_StdLogicVector(INIT_E)  &
                                                  To_StdLogicVector(INIT_D)  &
                                                  To_StdLogicVector(INIT_C)  &
                                                  To_StdLogicVector(INIT_B)  &
                                                  To_StdLogicVector(INIT_A)  &
                                                  To_StdLogicVector(INIT_9)  &
                                                  To_StdLogicVector(INIT_8)  &
                                                  To_StdLogicVector(INIT_7)  &
                                                  To_StdLogicVector(INIT_6)  &
                                                  To_StdLogicVector(INIT_5)  &
                                                  To_StdLogicVector(INIT_4)  &
                                                  To_StdLogicVector(INIT_3)  &
                                                  To_StdLogicVector(INIT_2)  &
                                                  To_StdLogicVector(INIT_1)  & 
                                                  To_StdLogicVector(INIT_0) ;  

  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLK'event and (WCLK = '1') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 1 loop
            MEM_temp(2*WADDR_in + i )  := WDATA(i) ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;


  end process ;


  ReadBehavior : process(RCLK)
  
    variable RADDR_in : integer range 0 to 8191 ;
    variable RDATA_temp : std_logic_vector( 1  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLK'event and (RCLK = '1') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 1 loop
            RDATA_temp(i ) := MEM(2*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;

  end process ;

end SB_RAM8192x2_ARCH;   --- SB_RAM8192x2


---------------------------------------
	--- SB_RAM8192x2NR
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM8192x2NR is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 1  downto 0) ;
                RCLKN : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'H';
                RADDR : in  std_logic_vector( 12  downto 0) ;
                WCLK  : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'H';
                WADDR : in  std_logic_vector( 12  downto 0) ;
                WDATA : in  std_logic_vector( 1  downto 0)
               );
  
  
end SB_RAM8192x2NR;

architecture SB_RAM8192x2NR_ARCH of SB_RAM8192x2NR is

  signal MEM : std_logic_vector(16383 downto 0) ;
  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLK)
    variable WADDR_in : integer range 0 to 8191;
    variable MEM_temp : std_logic_vector(16383 downto 0) :=  To_StdLogicVector(INIT_3F) &
                                                  To_StdLogicVector(INIT_3E) &
                                                  To_StdLogicVector(INIT_3D) &
                                                  To_StdLogicVector(INIT_3C) &
                                                  To_StdLogicVector(INIT_3B) &
                                                  To_StdLogicVector(INIT_3A) &
                                                  To_StdLogicVector(INIT_39) &
                                                  To_StdLogicVector(INIT_38) &
                                                  To_StdLogicVector(INIT_37) &
                                                  To_StdLogicVector(INIT_36) &
                                                  To_StdLogicVector(INIT_35) &
                                                  To_StdLogicVector(INIT_34) &
                                                  To_StdLogicVector(INIT_33) &
                                                  To_StdLogicVector(INIT_32) &
                                                  To_StdLogicVector(INIT_31) &
                                                  To_StdLogicVector(INIT_30) &
						  To_StdLogicVector(INIT_2F) &
                                                  To_StdLogicVector(INIT_2E) &
                                                  To_StdLogicVector(INIT_2D) &
                                                  To_StdLogicVector(INIT_2C) &
                                                  To_StdLogicVector(INIT_2B) &
                                                  To_StdLogicVector(INIT_2A) &
                                                  To_StdLogicVector(INIT_29) &
                                                  To_StdLogicVector(INIT_28) &
                                                  To_StdLogicVector(INIT_27) &
                                                  To_StdLogicVector(INIT_26) &
                                                  To_StdLogicVector(INIT_25) &
                                                  To_StdLogicVector(INIT_24) &
                                                  To_StdLogicVector(INIT_23) &
                                                  To_StdLogicVector(INIT_22) &
                                                  To_StdLogicVector(INIT_21) &
                                                  To_StdLogicVector(INIT_20) &
						  To_StdLogicVector(INIT_1F) &
                                                  To_StdLogicVector(INIT_1E) &
                                                  To_StdLogicVector(INIT_1D) &
                                                  To_StdLogicVector(INIT_1C) &
                                                  To_StdLogicVector(INIT_1B) &
                                                  To_StdLogicVector(INIT_1A) &
                                                  To_StdLogicVector(INIT_19) &
                                                  To_StdLogicVector(INIT_18) &
                                                  To_StdLogicVector(INIT_17) &
                                                  To_StdLogicVector(INIT_16) &
                                                  To_StdLogicVector(INIT_15) &
                                                  To_StdLogicVector(INIT_14) &
                                                  To_StdLogicVector(INIT_13) &
                                                  To_StdLogicVector(INIT_12) &
                                                  To_StdLogicVector(INIT_11) &
                                                  To_StdLogicVector(INIT_10) & 
						  To_StdLogicVector(INIT_F)  &
                                                  To_StdLogicVector(INIT_E)  &
                                                  To_StdLogicVector(INIT_D)  &
                                                  To_StdLogicVector(INIT_C)  &
                                                  To_StdLogicVector(INIT_B)  &
                                                  To_StdLogicVector(INIT_A)  &
                                                  To_StdLogicVector(INIT_9)  &
                                                  To_StdLogicVector(INIT_8)  &
                                                  To_StdLogicVector(INIT_7)  &
                                                  To_StdLogicVector(INIT_6)  &
                                                  To_StdLogicVector(INIT_5)  &
                                                  To_StdLogicVector(INIT_4)  &
                                                  To_StdLogicVector(INIT_3)  &
                                                  To_StdLogicVector(INIT_2)  &
                                                  To_StdLogicVector(INIT_1)  & 
                                                  To_StdLogicVector(INIT_0) ;  

  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLK'event and (WCLK = '1') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 1 loop
            MEM_temp(2*WADDR_in + i )  := WDATA(i) ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;


  end process ;


  ReadBehavior : process(RCLKN)
  
    variable RADDR_in : integer range 0 to 8191 ;
    variable RDATA_temp : std_logic_vector( 1  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLKN'event and (RCLKN = '0') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 1 loop
            RDATA_temp(i ) := MEM(2*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;

  end process ;

end SB_RAM8192x2NR_ARCH;   --- SB_RAM8192x2NR


---------------------------------------
	--- SB_RAM8192x2NW
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM8192x2NW is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 1  downto 0) ;
                RCLK  : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'H';
                RADDR : in  std_logic_vector( 12  downto 0) ;
                WCLKN : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'H';
                WADDR : in  std_logic_vector( 12  downto 0) ;
                WDATA : in  std_logic_vector( 1  downto 0)
               );
  
  
end SB_RAM8192x2NW;

architecture SB_RAM8192x2NW_ARCH of SB_RAM8192x2NW is
  
  signal MEM : std_logic_vector(16383 downto 0) ;
  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLKN)
    variable WADDR_in : integer range 0 to 8191;
    variable MEM_temp : std_logic_vector(16383 downto 0) :=  To_StdLogicVector(INIT_3F) &
                                                  To_StdLogicVector(INIT_3E) &
                                                  To_StdLogicVector(INIT_3D) &
                                                  To_StdLogicVector(INIT_3C) &
                                                  To_StdLogicVector(INIT_3B) &
                                                  To_StdLogicVector(INIT_3A) &
                                                  To_StdLogicVector(INIT_39) &
                                                  To_StdLogicVector(INIT_38) &
                                                  To_StdLogicVector(INIT_37) &
                                                  To_StdLogicVector(INIT_36) &
                                                  To_StdLogicVector(INIT_35) &
                                                  To_StdLogicVector(INIT_34) &
                                                  To_StdLogicVector(INIT_33) &
                                                  To_StdLogicVector(INIT_32) &
                                                  To_StdLogicVector(INIT_31) &
                                                  To_StdLogicVector(INIT_30) &
						  To_StdLogicVector(INIT_2F) &
                                                  To_StdLogicVector(INIT_2E) &
                                                  To_StdLogicVector(INIT_2D) &
                                                  To_StdLogicVector(INIT_2C) &
                                                  To_StdLogicVector(INIT_2B) &
                                                  To_StdLogicVector(INIT_2A) &
                                                  To_StdLogicVector(INIT_29) &
                                                  To_StdLogicVector(INIT_28) &
                                                  To_StdLogicVector(INIT_27) &
                                                  To_StdLogicVector(INIT_26) &
                                                  To_StdLogicVector(INIT_25) &
                                                  To_StdLogicVector(INIT_24) &
                                                  To_StdLogicVector(INIT_23) &
                                                  To_StdLogicVector(INIT_22) &
                                                  To_StdLogicVector(INIT_21) &
                                                  To_StdLogicVector(INIT_20) &
						  To_StdLogicVector(INIT_1F) &
                                                  To_StdLogicVector(INIT_1E) &
                                                  To_StdLogicVector(INIT_1D) &
                                                  To_StdLogicVector(INIT_1C) &
                                                  To_StdLogicVector(INIT_1B) &
                                                  To_StdLogicVector(INIT_1A) &
                                                  To_StdLogicVector(INIT_19) &
                                                  To_StdLogicVector(INIT_18) &
                                                  To_StdLogicVector(INIT_17) &
                                                  To_StdLogicVector(INIT_16) &
                                                  To_StdLogicVector(INIT_15) &
                                                  To_StdLogicVector(INIT_14) &
                                                  To_StdLogicVector(INIT_13) &
                                                  To_StdLogicVector(INIT_12) &
                                                  To_StdLogicVector(INIT_11) &
                                                  To_StdLogicVector(INIT_10) & 
						  To_StdLogicVector(INIT_F)  &
                                                  To_StdLogicVector(INIT_E)  &
                                                  To_StdLogicVector(INIT_D)  &
                                                  To_StdLogicVector(INIT_C)  &
                                                  To_StdLogicVector(INIT_B)  &
                                                  To_StdLogicVector(INIT_A)  &
                                                  To_StdLogicVector(INIT_9)  &
                                                  To_StdLogicVector(INIT_8)  &
                                                  To_StdLogicVector(INIT_7)  &
                                                  To_StdLogicVector(INIT_6)  &
                                                  To_StdLogicVector(INIT_5)  &
                                                  To_StdLogicVector(INIT_4)  &
                                                  To_StdLogicVector(INIT_3)  &
                                                  To_StdLogicVector(INIT_2)  &
                                                  To_StdLogicVector(INIT_1)  & 
                                                  To_StdLogicVector(INIT_0) ;  

  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLKN'event and (WCLKN = '0') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 1 loop
            MEM_temp(2*WADDR_in + i )  := WDATA(i) ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;


  end process ;


  ReadBehavior : process(RCLK)
  
    variable RADDR_in : integer range 0 to 8191 ;
    variable RDATA_temp : std_logic_vector( 1  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLK'event and (RCLK = '1') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 1 loop
            RDATA_temp(i ) := MEM(2*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;

  end process ;

end SB_RAM8192x2NW_ARCH;   --- SB_RAM8192x2NW


---------------------------------------
	--- SB_RAM8192x2NRNW
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM8192x2NRNW is

  generic ( 
           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 1  downto 0) ;
                RCLKN : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'H';
                RADDR : in  std_logic_vector( 12  downto 0) ;
                WCLKN : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'H';
                WADDR : in  std_logic_vector( 12  downto 0) ;
                WDATA : in  std_logic_vector( 1  downto 0)
               );
  
  
end SB_RAM8192x2NRNW;

architecture SB_RAM8192x2NRNW_ARCH of SB_RAM8192x2NRNW is
 
  signal MEM : std_logic_vector(16383 downto 0) ;
  signal Address_Collision_Detected : std_logic ;

begin 

  process(RE,WE,WADDR,RADDR)
      begin
          if ( (WE = '1')  and (RE = '1') and ( WADDR = RADDR) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;

          assert (Address_Collision_Detected = '0')
            report "Address_Collision"
            severity warning ; 
  end process; 

  WriteBehavior : process(WCLKN)
    variable WADDR_in : integer range 0 to 8191;
    variable MEM_temp : std_logic_vector(16383 downto 0) :=  To_StdLogicVector(INIT_3F) &
                                                  To_StdLogicVector(INIT_3E) &
                                                  To_StdLogicVector(INIT_3D) &
                                                  To_StdLogicVector(INIT_3C) &
                                                  To_StdLogicVector(INIT_3B) &
                                                  To_StdLogicVector(INIT_3A) &
                                                  To_StdLogicVector(INIT_39) &
                                                  To_StdLogicVector(INIT_38) &
                                                  To_StdLogicVector(INIT_37) &
                                                  To_StdLogicVector(INIT_36) &
                                                  To_StdLogicVector(INIT_35) &
                                                  To_StdLogicVector(INIT_34) &
                                                  To_StdLogicVector(INIT_33) &
                                                  To_StdLogicVector(INIT_32) &
                                                  To_StdLogicVector(INIT_31) &
                                                  To_StdLogicVector(INIT_30) &
						  To_StdLogicVector(INIT_2F) &
                                                  To_StdLogicVector(INIT_2E) &
                                                  To_StdLogicVector(INIT_2D) &
                                                  To_StdLogicVector(INIT_2C) &
                                                  To_StdLogicVector(INIT_2B) &
                                                  To_StdLogicVector(INIT_2A) &
                                                  To_StdLogicVector(INIT_29) &
                                                  To_StdLogicVector(INIT_28) &
                                                  To_StdLogicVector(INIT_27) &
                                                  To_StdLogicVector(INIT_26) &
                                                  To_StdLogicVector(INIT_25) &
                                                  To_StdLogicVector(INIT_24) &
                                                  To_StdLogicVector(INIT_23) &
                                                  To_StdLogicVector(INIT_22) &
                                                  To_StdLogicVector(INIT_21) &
                                                  To_StdLogicVector(INIT_20) &
						  To_StdLogicVector(INIT_1F) &
                                                  To_StdLogicVector(INIT_1E) &
                                                  To_StdLogicVector(INIT_1D) &
                                                  To_StdLogicVector(INIT_1C) &
                                                  To_StdLogicVector(INIT_1B) &
                                                  To_StdLogicVector(INIT_1A) &
                                                  To_StdLogicVector(INIT_19) &
                                                  To_StdLogicVector(INIT_18) &
                                                  To_StdLogicVector(INIT_17) &
                                                  To_StdLogicVector(INIT_16) &
                                                  To_StdLogicVector(INIT_15) &
                                                  To_StdLogicVector(INIT_14) &
                                                  To_StdLogicVector(INIT_13) &
                                                  To_StdLogicVector(INIT_12) &
                                                  To_StdLogicVector(INIT_11) &
                                                  To_StdLogicVector(INIT_10) & 
						  To_StdLogicVector(INIT_F)  &
                                                  To_StdLogicVector(INIT_E)  &
                                                  To_StdLogicVector(INIT_D)  &
                                                  To_StdLogicVector(INIT_C)  &
                                                  To_StdLogicVector(INIT_B)  &
                                                  To_StdLogicVector(INIT_A)  &
                                                  To_StdLogicVector(INIT_9)  &
                                                  To_StdLogicVector(INIT_8)  &
                                                  To_StdLogicVector(INIT_7)  &
                                                  To_StdLogicVector(INIT_6)  &
                                                  To_StdLogicVector(INIT_5)  &
                                                  To_StdLogicVector(INIT_4)  &
                                                  To_StdLogicVector(INIT_3)  &
                                                  To_StdLogicVector(INIT_2)  &
                                                  To_StdLogicVector(INIT_1)  & 
                                                  To_StdLogicVector(INIT_0) ;  

  begin

    WADDR_in := conv_integer(WADDR) ;
  
    if ( WCLKN'event and (WCLKN = '0') and (WCLKE = '1') and (WE = '1') ) then
       for i in 0 to 1 loop
            MEM_temp(2*WADDR_in + i )  := WDATA(i) ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;


  end process ;


  ReadBehavior : process(RCLKN)
  
    variable RADDR_in : integer range 0 to 8191 ;
    variable RDATA_temp : std_logic_vector( 1  downto 0) ; 
    
  begin 

    RADDR_in := conv_integer(RADDR) ;

    if ( Address_Collision_Detected = '1') then
        RDATA_temp := (others => 'X') ;
    elsif ( RCLKN'event and (RCLKN = '0') and (RCLKE = '1') and (RE = '1') ) then
       for i in 0 to 1 loop
            RDATA_temp(i ) := MEM(2*RADDR_in + i )  ;
       end loop ;
    end if ; 

    RDATA <= RDATA_temp ;

  end process ;
end SB_RAM8192x2NRNW_ARCH;   --- SB_RAM8192x2NRNW

-------------------------------------------------------------------
--    SB_RAM16K Leaf Level Ram Block for 16K Physical Ram Wrappers   
-------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
use IEEE.VITAL_Timing.all; 
USE IEEE.numeric_std.ALL;

entity SB_RAM16K is

  generic ( 
           TimingChecksOn : boolean := true;
           Xon            : boolean := false;
           MsgOn          : boolean := false;
           
           tipd_RCLK  : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_RCLKE : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_RE    : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_RADDR : VitalDelayArrayType01(9 downto 0)  := (others => (0 ns, 0 ns));
           tipd_WCLK  : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_WCLKE : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_WE    : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_WADDR : VitalDelayArrayType01(9 downto 0)  := (others => (0 ns, 0 ns));
           tipd_MASK  : VitalDelayArrayType01(15 downto 0)  := (others => (0 ns, 0 ns));
           tipd_WDATA : VitalDelayArrayType01(15 downto 0)  := (others => (0 ns, 0 ns));

           tpd_RCLK_RDATA : VitalDelayArrayType01(15 downto 0) := (others => (100 ns, 100 ns));
           tpd_RCLK_RDATA_posedge : VitalDelayArrayType01(15 downto 0) := (others => (100 ns, 100 ns));

           tsetup_RADDR_RCLK_negedge_posedge : VitalDelayArrayType(9 downto 0)  := (others => 0 ns);
           tsetup_RADDR_RCLK_posedge_posedge : VitalDelayArrayType(9 downto 0)  := (others => 0 ns);
           tsetup_RCLKE_RCLK_negedge_posedge : VitalDelayType                   := 0 ns;
           tsetup_RCLKE_RCLK_posedge_posedge : VitalDelayType                   := 0 ns;
           tsetup_RE_RCLK_negedge_posedge    : VitalDelayType                   := 0 ns;
           tsetup_RE_RCLK_posedge_posedge    : VitalDelayType                   := 0 ns;

           tsetup_WADDR_WCLK_negedge_posedge : VitalDelayArrayType(9 downto 0)  := (others => 0 ns);
           tsetup_WADDR_WCLK_posedge_posedge : VitalDelayArrayType(9 downto 0)  := (others => 0 ns);
           tsetup_WDATA_WCLK_negedge_posedge : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           tsetup_WDATA_WCLK_posedge_posedge : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           tsetup_WCLKE_WCLK_negedge_posedge : VitalDelayType                   := 0 ns;
           tsetup_WCLKE_WCLK_posedge_posedge : VitalDelayType                   := 0 ns;
           tsetup_WE_WCLK_negedge_posedge    : VitalDelayType                   := 0 ns;
           tsetup_WE_WCLK_posedge_posedge    : VitalDelayType                   := 0 ns;
           tsetup_MASK_WCLK_negedge_posedge  : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           tsetup_MASK_WCLK_posedge_posedge  : VitalDelayArrayType(15 downto 0) := (others => 0 ns);

           thold_RADDR_RCLK_negedge_posedge : VitalDelayArrayType(9 downto 0)  := (others => 0 ns);
           thold_RADDR_RCLK_posedge_posedge : VitalDelayArrayType(9 downto 0)  := (others => 0 ns);
           thold_RCLKE_RCLK_negedge_posedge : VitalDelayType                   := 0 ns;
           thold_RCLKE_RCLK_posedge_posedge : VitalDelayType                   := 0 ns;
           thold_RE_RCLK_negedge_posedge    : VitalDelayType                   := 0 ns;
           thold_RE_RCLK_posedge_posedge    : VitalDelayType                   := 0 ns;

           thold_WADDR_WCLK_negedge_posedge : VitalDelayArrayType(9 downto 0)  := (others => 0 ns);
           thold_WADDR_WCLK_posedge_posedge : VitalDelayArrayType(9 downto 0)  := (others => 0 ns);
           thold_WDATA_WCLK_negedge_posedge : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           thold_WDATA_WCLK_posedge_posedge : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           thold_WCLKE_WCLK_negedge_posedge : VitalDelayType                   := 0 ns;
           thold_WCLKE_WCLK_posedge_posedge : VitalDelayType                   := 0 ns;
           thold_WE_WCLK_negedge_posedge    : VitalDelayType                   := 0 ns;
           thold_WE_WCLK_posedge_posedge    : VitalDelayType                   := 0 ns;
           thold_MASK_WCLK_negedge_posedge  : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           thold_MASK_WCLK_posedge_posedge  : VitalDelayArrayType(15 downto 0) := (others => 0 ns);

           tpw_RCLK_negedge : VitalDelayType := 0 ns;
           tpw_RCLK_posedge : VitalDelayType := 0 ns;
           tpw_WCLK_negedge : VitalDelayType := 0 ns;
           tpw_WCLK_posedge : VitalDelayType := 0 ns;


           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
 
           INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 15  downto 0) ;
                RCLK  : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'L';
                RADDR : in  std_logic_vector( 9  downto 0) ;
                WCLK  : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'L';
                WADDR : in  std_logic_vector( 9  downto 0) ;
                MASK  : in  std_logic_vector( 15  downto 0) ;
                WDATA : in  std_logic_vector( 15  downto 0)
               );
  
end SB_RAM16K;



architecture SB_RAM16K_V of SB_RAM16K is

  signal MEM : std_logic_vector(16383 downto 0) ;
  signal Address_Collision_Detected : std_logic ;


  signal RADDR_ipd : std_logic_vector(9 downto 0)  := (others => 'X');   
  signal RCLK_ipd  : std_logic                    := 'X';
  signal RCLKE_ipd : std_logic                    := 'X';
  signal RE_ipd    : std_logic                    := 'X';

  signal WADDR_ipd : std_logic_vector(9 downto 0)  := (others => 'X');
  signal WCLK_ipd  : std_logic                    := 'X';  
  signal WCLKE_ipd : std_logic                    := 'X';
  signal WE_ipd    : std_logic                    := 'X';
  signal MASK_ipd  : std_logic_vector(15 downto 0) := (others => 'X');
  signal WDATA_ipd : std_logic_vector(15 downto 0) := (others => 'X');

  signal RADDR_in : integer range 0 to 1023;  -- 1Kx16 
  signal WADDR_in : integer range 0 to 1023; 

begin

---------------------
--  Input Wire Delay
---------------------
  WireDelay : block
  begin
    RADDR_DELAY : for i in 9 downto 0 generate
       VitalWireDelay (RADDR_ipd(i), RADDR(i), tipd_RADDR(i));
    end generate RADDR_DELAY;
    VitalWireDelay (RCLK_ipd, RCLK, tipd_RCLK);
    VitalWireDelay (RCLKE_ipd, RCLKE, tipd_RCLKE);
    VitalWireDelay (RE_ipd, RE, tipd_RE);
    WADDR_DELAY : for i in 9 downto 0 generate
       VitalWireDelay (WADDR_ipd(i), WADDR(i), tipd_WADDR(i));
    end generate WADDR_DELAY;
    VitalWireDelay (WCLK_ipd, WCLK, tipd_WCLK);
    VitalWireDelay (WCLKE_ipd, WCLKE, tipd_WCLKE);
    VitalWireDelay (WE_ipd, WE, tipd_WE);
    MASK_DELAY : for i in 15 downto 0 generate
       VitalWireDelay (MASK_ipd(i), MASK(i), tipd_MASK(i));
    end generate MASK_DELAY;
    WDATA_DELAY : for i in 15 downto 0 generate
       VitalWireDelay (WDATA_ipd(i), WDATA(i), tipd_WDATA(i));
    end generate WDATA_DELAY;
  end block;

  process(RE_ipd,WE_ipd,WADDR_ipd,RADDR_ipd)
      begin
          if ( (WE_ipd = '1')  and (RE_ipd = '1') and ( WADDR_ipd = RADDR_ipd) ) then
             Address_Collision_Detected <= '1';
          else
             Address_Collision_Detected <= '0' ;
          end if ;
          assert (not(Address_Collision_Detected = '1'))
            report "Address_Collision"
            severity warning ;         
  end process; 



  VITALReadBehavior : process(RADDR_ipd,RCLK_ipd,RCLKE_ipd,RE_ipd)
   
       variable Tviol_RADDR0_RCLK_posedge : std_logic := '0';
       variable Tviol_RADDR1_RCLK_posedge : std_logic := '0';
       variable Tviol_RADDR2_RCLK_posedge : std_logic := '0';
       variable Tviol_RADDR3_RCLK_posedge : std_logic := '0';
       variable Tviol_RADDR4_RCLK_posedge : std_logic := '0';
       variable Tviol_RADDR5_RCLK_posedge : std_logic := '0';
       variable Tviol_RADDR6_RCLK_posedge : std_logic := '0';
       variable Tviol_RADDR7_RCLK_posedge : std_logic := '0';
       variable Tviol_RADDR8_RCLK_posedge : std_logic := '0';
       variable Tviol_RADDR9_RCLK_posedge : std_logic := '0';
       variable Tviol_RCLKE_RCLK_posedge  : std_logic := '0';
       variable Tviol_RE_RCLK_posedge     : std_logic := '0';

       variable Tmkr_RADDR0_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR1_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR2_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR3_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR4_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR5_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR6_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR7_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR8_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RADDR9_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RCLKE_RCLK_posedge  : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_RE_RCLK_posedge     : VitalTimingDataType := VitalTimingDataInit;

       variable PViol_RCLK : std_logic := '0';

       variable PInfo_RCLK : VitalPeriodDataType ;

       variable RDATA_GlitchData0  : VitalGlitchDataType;
       variable RDATA_GlitchData1  : VitalGlitchDataType;
       variable RDATA_GlitchData2  : VitalGlitchDataType;
       variable RDATA_GlitchData3  : VitalGlitchDataType;
       variable RDATA_GlitchData4  : VitalGlitchDataType;
       variable RDATA_GlitchData5  : VitalGlitchDataType;
       variable RDATA_GlitchData6  : VitalGlitchDataType;
       variable RDATA_GlitchData7  : VitalGlitchDataType;
       variable RDATA_GlitchData8  : VitalGlitchDataType;
       variable RDATA_GlitchData9  : VitalGlitchDataType;
       variable RDATA_GlitchData10 : VitalGlitchDataType;
       variable RDATA_GlitchData11 : VitalGlitchDataType;
       variable RDATA_GlitchData12 : VitalGlitchDataType;
       variable RDATA_GlitchData13 : VitalGlitchDataType;
       variable RDATA_GlitchData14 : VitalGlitchDataType;
       variable RDATA_GlitchData15 : VitalGlitchDataType;

       variable Violation     : std_logic  := '0';

       variable temp : std_logic_vector(15 downto 0) := (others => 'X');   --X 
       variable RDATA_zd : std_logic_vector(15 downto 0) := (others => 'X'); --X 

  begin

  -------------------------
  --  Functionality Section
  -------------------------
    RADDR_in <= conv_integer(RADDR_ipd) ;
  
    if (Violation = '1') then
       RDATA <= (others => 'X') ;
    elsif ( RCLK_ipd'event and (RCLK_ipd = '1') and (RCLKE_ipd = '1' or RCLKE_ipd = 'H') and (RE_ipd = '1') ) then
       for i in 0 to 15 loop
         temp(i) := MEM(16*RADDR_in + i ) ;
       end loop ;
    end if ; 

    RDATA <= temp;


  ------------------------
  --  Timing Check Section
  ------------------------
    if (TimingChecksOn) then
      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR0_RCLK_posedge,
        TimingData     => Tmkr_RADDR0_RCLK_posedge,
        TestSignal     => RADDR_ipd(0),
        TestSignalName => "RADDR(0)",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(0),
        SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(0),
        HoldLow        => thold_RADDR_RCLK_posedge_posedge(0),
        HoldHigh       => thold_RADDR_RCLK_negedge_posedge(0),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR1_RCLK_posedge,
        TimingData     => Tmkr_RADDR1_RCLK_posedge,
        TestSignal     => RADDR_ipd(1),
        TestSignalName => "RADDR(1)",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(1),
        SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(1),
        HoldLow        => thold_RADDR_RCLK_posedge_posedge(1),
        HoldHigh       => thold_RADDR_RCLK_negedge_posedge(1),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR2_RCLK_posedge,
        TimingData     => Tmkr_RADDR2_RCLK_posedge,
        TestSignal     => RADDR_ipd(2),
        TestSignalName => "RADDR(2)",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(2),
        SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(2),
        HoldLow        => thold_RADDR_RCLK_posedge_posedge(2),
        HoldHigh       => thold_RADDR_RCLK_negedge_posedge(2),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR3_RCLK_posedge,
        TimingData     => Tmkr_RADDR3_RCLK_posedge,
        TestSignal     => RADDR_ipd(3),
        TestSignalName => "RADDR(3)",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(3),
        SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(3),
        HoldLow        => thold_RADDR_RCLK_posedge_posedge(3),
        HoldHigh       => thold_RADDR_RCLK_negedge_posedge(3),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR4_RCLK_posedge,
        TimingData     => Tmkr_RADDR4_RCLK_posedge,
        TestSignal     => RADDR_ipd(4),
        TestSignalName => "RADDR(4)",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(4),
        SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(4),
        HoldLow        => thold_RADDR_RCLK_posedge_posedge(4),
        HoldHigh       => thold_RADDR_RCLK_negedge_posedge(4),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR5_RCLK_posedge,
        TimingData     => Tmkr_RADDR5_RCLK_posedge,
        TestSignal     => RADDR_ipd(5),
        TestSignalName => "RADDR(5)",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(5),
        SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(5),
        HoldLow        => thold_RADDR_RCLK_posedge_posedge(5),
        HoldHigh       => thold_RADDR_RCLK_negedge_posedge(5),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR6_RCLK_posedge,
        TimingData     => Tmkr_RADDR6_RCLK_posedge,
        TestSignal     => RADDR_ipd(6),
        TestSignalName => "RADDR(6)",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(6),
        SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(6),
        HoldLow        => thold_RADDR_RCLK_posedge_posedge(6),
        HoldHigh       => thold_RADDR_RCLK_negedge_posedge(6),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR7_RCLK_posedge,
        TimingData     => Tmkr_RADDR7_RCLK_posedge,
        TestSignal     => RADDR_ipd(7),
        TestSignalName => "RADDR(7)",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(7),
        SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(7),
        HoldLow        => thold_RADDR_RCLK_posedge_posedge(7),
        HoldHigh       => thold_RADDR_RCLK_negedge_posedge(7),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);


      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR8_RCLK_posedge,
        TimingData     => Tmkr_RADDR8_RCLK_posedge,
        TestSignal     => RADDR_ipd(8),
        TestSignalName => "RADDR(8)",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(8),
        SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(8),
        HoldLow        => thold_RADDR_RCLK_posedge_posedge(8),
        HoldHigh       => thold_RADDR_RCLK_negedge_posedge(8),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);


      VitalSetupHoldCheck (
        Violation      => Tviol_RADDR9_RCLK_posedge,
        TimingData     => Tmkr_RADDR9_RCLK_posedge,
        TestSignal     => RADDR_ipd(9),
        TestSignalName => "RADDR(9)",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(9),
        SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(9),
        HoldLow        => thold_RADDR_RCLK_posedge_posedge(9),
        HoldHigh       => thold_RADDR_RCLK_negedge_posedge(9),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_RCLKE_RCLK_posedge,
        TimingData     => Tmkr_RCLKE_RCLK_posedge,
        TestSignal     => RCLKE_ipd,
        TestSignalName => "RCLKE",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RCLKE_RCLK_posedge_posedge,
        SetupLow       => tsetup_RCLKE_RCLK_negedge_posedge,
        HoldLow        => thold_RCLKE_RCLK_posedge_posedge,
        HoldHigh       => thold_RCLKE_RCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_RE_RCLK_posedge,
        TimingData     => Tmkr_RE_RCLK_posedge,
        TestSignal     => RCLK_ipd,
        TestSignalName => "RCLK",
        TestDelay      => 0 ns,
        RefSignal      => RCLK_ipd,
        RefSignalName  => "RCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_RE_RCLK_posedge_posedge,
        SetupLow       => tsetup_RE_RCLK_negedge_posedge,
        HoldLow        => thold_RE_RCLK_posedge_posedge,
        HoldHigh       => thold_RE_RCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
               

      VitalPeriodPulseCheck (
        Violation      => Pviol_RCLK,
        PeriodData     => PInfo_RCLK,
        TestSignal     => RCLK_ipd,
        TestSignalName => "RCLK",
        TestDelay      => 0 ns,
        Period         => 0 ns,
        PulseWidthHigh => tpw_RCLK_posedge,
        PulseWidthLow  => tpw_RCLK_negedge,
        CheckEnabled   => true,
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

    end if ;

    Violation  := Pviol_RCLK or
                  Tviol_RADDR0_RCLK_posedge or
                  Tviol_RADDR1_RCLK_posedge or
                  Tviol_RADDR2_RCLK_posedge or
                  Tviol_RADDR3_RCLK_posedge or
                  Tviol_RADDR4_RCLK_posedge or
                  Tviol_RADDR5_RCLK_posedge or
                  Tviol_RADDR6_RCLK_posedge or
                  Tviol_RADDR7_RCLK_posedge or
                  Tviol_RCLKE_RCLK_posedge or
                  Tviol_RE_RCLK_posedge;

    RDATA_zd(0) := Violation xor RDATA_zd(0) ;
    RDATA_zd(1) := Violation xor RDATA_zd(1) ;
    RDATA_zd(2) := Violation xor RDATA_zd(2) ;
    RDATA_zd(3) := Violation xor RDATA_zd(3) ;
    RDATA_zd(4) := Violation xor RDATA_zd(4) ;
    RDATA_zd(5) := Violation xor RDATA_zd(5) ;
    RDATA_zd(6) := Violation xor RDATA_zd(6) ;
    RDATA_zd(7) := Violation xor RDATA_zd(7) ;
    RDATA_zd(8) := Violation xor RDATA_zd(8) ;
    RDATA_zd(9) := Violation xor RDATA_zd(9) ;
    RDATA_zd(10) := Violation xor RDATA_zd(10) ;
    RDATA_zd(11) := Violation xor RDATA_zd(11) ;
    RDATA_zd(12) := Violation xor RDATA_zd(12) ;
    RDATA_zd(13) := Violation xor RDATA_zd(13) ;
    RDATA_zd(14) := Violation xor RDATA_zd(14) ;
    RDATA_zd(15) := Violation xor RDATA_zd(15) ;
    
    
  ----------------------
  --  Path Delay Section
  ----------------------
    VitalPathDelay01 (
      OutSignal     => RDATA(0),
      GlitchData    => RDATA_GlitchData0,
      OutSignalName => "RDATA(0)",
      OutTemp       => RDATA_zd(0),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(0), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(1),
      GlitchData    => RDATA_GlitchData1,
      OutSignalName => "RDATA(1)",
      OutTemp       => RDATA_zd(1),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(1), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(2),
      GlitchData    => RDATA_GlitchData2,
      OutSignalName => "RDATA(2)",
      OutTemp       => RDATA_zd(2),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(2), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(3),
      GlitchData    => RDATA_GlitchData3,
      OutSignalName => "RDATA(3)",
      OutTemp       => RDATA_zd(3),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(3), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(4),
      GlitchData    => RDATA_GlitchData4,
      OutSignalName => "RDATA(4)",
      OutTemp       => RDATA_zd(4),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(4), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(5),
      GlitchData    => RDATA_GlitchData5,
      OutSignalName => "RDATA(5)",
      OutTemp       => RDATA_zd(5),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(5), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(6),
      GlitchData    => RDATA_GlitchData6,
      OutSignalName => "RDATA(6)",
      OutTemp       => RDATA_zd(6),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(6), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(7),
      GlitchData    => RDATA_GlitchData7,
      OutSignalName => "RDATA(7)",
      OutTemp       => RDATA_zd(7),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(7), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(8),
      GlitchData    => RDATA_GlitchData8,
      OutSignalName => "RDATA(8)",
      OutTemp       => RDATA_zd(8),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(8), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(9),
      GlitchData    => RDATA_GlitchData9,
      OutSignalName => "RDATA(9)",
      OutTemp       => RDATA_zd(9),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(9), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(10),
      GlitchData    => RDATA_GlitchData10,
      OutSignalName => "RDATA(10)",
      OutTemp       => RDATA_zd(10),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(10), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(11),
      GlitchData    => RDATA_GlitchData11,
      OutSignalName => "RDATA(11)",
      OutTemp       => RDATA_zd(11),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(11), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(12),
      GlitchData    => RDATA_GlitchData12,
      OutSignalName => "RDATA(12)",
      OutTemp       => RDATA_zd(12),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(12), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(13),
      GlitchData    => RDATA_GlitchData13,
      OutSignalName => "RDATA(13)",
      OutTemp       => RDATA_zd(13),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(13), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(14),
      GlitchData    => RDATA_GlitchData14,
      OutSignalName => "RDATA(14)",
      OutTemp       => RDATA_zd(14),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(14), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(15),
      GlitchData    => RDATA_GlitchData15,
      OutSignalName => "RDATA(15)",
      OutTemp       => RDATA_zd(15),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(15), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(0),
      GlitchData    => RDATA_GlitchData0,
      OutSignalName => "RDATA(0)",
      OutTemp       => RDATA_zd(0),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(0), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(1),
      GlitchData    => RDATA_GlitchData1,
      OutSignalName => "RDATA(1)",
      OutTemp       => RDATA_zd(1),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(1), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(2),
      GlitchData    => RDATA_GlitchData2,
      OutSignalName => "RDATA(2)",
      OutTemp       => RDATA_zd(2),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(2), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(3),
      GlitchData    => RDATA_GlitchData3,
      OutSignalName => "RDATA(3)",
      OutTemp       => RDATA_zd(3),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(3), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(4),
      GlitchData    => RDATA_GlitchData4,
      OutSignalName => "RDATA(4)",
      OutTemp       => RDATA_zd(4),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(4), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(5),
      GlitchData    => RDATA_GlitchData5,
      OutSignalName => "RDATA(5)",
      OutTemp       => RDATA_zd(5),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(5), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(6),
      GlitchData    => RDATA_GlitchData6,
      OutSignalName => "RDATA(6)",
      OutTemp       => RDATA_zd(6),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(6), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(7),
      GlitchData    => RDATA_GlitchData7,
      OutSignalName => "RDATA(7)",
      OutTemp       => RDATA_zd(7),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(7), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(8),
      GlitchData    => RDATA_GlitchData8,
      OutSignalName => "RDATA(8)",
      OutTemp       => RDATA_zd(8),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(8), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(9),
      GlitchData    => RDATA_GlitchData9,
      OutSignalName => "RDATA(9)",
      OutTemp       => RDATA_zd(9),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(9), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(10),
      GlitchData    => RDATA_GlitchData10,
      OutSignalName => "RDATA(10)",
      OutTemp       => RDATA_zd(10),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(10), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(11),
      GlitchData    => RDATA_GlitchData11,
      OutSignalName => "RDATA(11)",
      OutTemp       => RDATA_zd(11),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(11), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(12),
      GlitchData    => RDATA_GlitchData12,
      OutSignalName => "RDATA(12)",
      OutTemp       => RDATA_zd(12),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(12), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(13),
      GlitchData    => RDATA_GlitchData13,
      OutSignalName => "RDATA(13)",
      OutTemp       => RDATA_zd(13),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(13), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(14),
      GlitchData    => RDATA_GlitchData14,
      OutSignalName => "RDATA(14)",
      OutTemp       => RDATA_zd(14),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(14), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

    VitalPathDelay01 (
      OutSignal     => RDATA(15),
      GlitchData    => RDATA_GlitchData15,
      OutSignalName => "RDATA(15)",
      OutTemp       => RDATA_zd(15),
      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA_posedge(15), true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);

  end process VITALReadBehavior;



  VITALWriteBehavior : process(WADDR_ipd,WCLK_ipd,WCLKE_ipd,WE_ipd,MASK_ipd) 

       variable Tviol_WADDR0_WCLK_posedge : std_logic := '0';
       variable Tviol_WADDR1_WCLK_posedge : std_logic := '0';
       variable Tviol_WADDR2_WCLK_posedge : std_logic := '0';
       variable Tviol_WADDR3_WCLK_posedge : std_logic := '0';
       variable Tviol_WADDR4_WCLK_posedge : std_logic := '0';
       variable Tviol_WADDR5_WCLK_posedge : std_logic := '0';
       variable Tviol_WADDR6_WCLK_posedge : std_logic := '0';
       variable Tviol_WADDR7_WCLK_posedge : std_logic := '0';
       variable Tviol_WADDR8_WCLK_posedge : std_logic := '0';
       variable Tviol_WADDR9_WCLK_posedge : std_logic := '0';
       variable Tviol_WCLKE_WCLK_posedge  : std_logic := '0';
       variable Tviol_WE_WCLK_posedge     : std_logic := '0';
       variable Tviol_WDATA0_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA1_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA2_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA3_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA4_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA5_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA6_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA7_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA8_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA9_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA10_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA11_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA12_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA13_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA14_WCLK_posedge : std_logic := '0';
       variable Tviol_WDATA15_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK0_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK1_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK2_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK3_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK4_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK5_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK6_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK7_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK8_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK9_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK10_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK11_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK12_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK13_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK14_WCLK_posedge : std_logic := '0';
       variable Tviol_MASK15_WCLK_posedge : std_logic := '0';


       variable Tmkr_WADDR0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR5_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR6_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR7_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR8_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WADDR9_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WCLKE_WCLK_posedge  : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WE_WCLK_posedge     : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA5_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA6_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA7_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA8_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA9_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA10_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA11_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA12_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA13_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA14_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_WDATA15_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK5_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK6_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK7_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK8_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK9_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK10_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK11_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK12_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK13_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK14_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
       variable Tmkr_MASK15_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;

       variable PViol_WCLK : std_logic := '0';

       variable PInfo_WCLK : VitalPeriodDataType := VitalPeriodDataInit;


       variable Violation     : std_logic  := '0';
       variable MEM_temp : std_logic_vector(16383 downto 0) :=  To_StdLogicVector(INIT_3F) &
                                                  To_StdLogicVector(INIT_3E) &
                                                  To_StdLogicVector(INIT_3D) &
                                                  To_StdLogicVector(INIT_3C) &
                                                  To_StdLogicVector(INIT_3B) &
                                                  To_StdLogicVector(INIT_3A) &
                                                  To_StdLogicVector(INIT_39) &
                                                  To_StdLogicVector(INIT_38) &
                                                  To_StdLogicVector(INIT_37) &
                                                  To_StdLogicVector(INIT_36) &
                                                  To_StdLogicVector(INIT_35) &
                                                  To_StdLogicVector(INIT_34) &
                                                  To_StdLogicVector(INIT_33) &
                                                  To_StdLogicVector(INIT_32) &
                                                  To_StdLogicVector(INIT_31) &
                                                  To_StdLogicVector(INIT_30) &
						  To_StdLogicVector(INIT_2F) &
                                                  To_StdLogicVector(INIT_2E) &
                                                  To_StdLogicVector(INIT_2D) &
                                                  To_StdLogicVector(INIT_2C) &
                                                  To_StdLogicVector(INIT_2B) &
                                                  To_StdLogicVector(INIT_2A) &
                                                  To_StdLogicVector(INIT_29) &
                                                  To_StdLogicVector(INIT_28) &
                                                  To_StdLogicVector(INIT_27) &
                                                  To_StdLogicVector(INIT_26) &
                                                  To_StdLogicVector(INIT_25) &
                                                  To_StdLogicVector(INIT_24) &
                                                  To_StdLogicVector(INIT_23) &
                                                  To_StdLogicVector(INIT_22) &
                                                  To_StdLogicVector(INIT_21) &
                                                  To_StdLogicVector(INIT_20) &
						  To_StdLogicVector(INIT_1F) &
                                                  To_StdLogicVector(INIT_1E) &
                                                  To_StdLogicVector(INIT_1D) &
                                                  To_StdLogicVector(INIT_1C) &
                                                  To_StdLogicVector(INIT_1B) &
                                                  To_StdLogicVector(INIT_1A) &
                                                  To_StdLogicVector(INIT_19) &
                                                  To_StdLogicVector(INIT_18) &
                                                  To_StdLogicVector(INIT_17) &
                                                  To_StdLogicVector(INIT_16) &
                                                  To_StdLogicVector(INIT_15) &
                                                  To_StdLogicVector(INIT_14) &
                                                  To_StdLogicVector(INIT_13) &
                                                  To_StdLogicVector(INIT_12) &
                                                  To_StdLogicVector(INIT_11) &
                                                  To_StdLogicVector(INIT_10) & 
						  To_StdLogicVector(INIT_F)  &
                                                  To_StdLogicVector(INIT_E)  &
                                                  To_StdLogicVector(INIT_D)  &
                                                  To_StdLogicVector(INIT_C)  &
                                                  To_StdLogicVector(INIT_B)  &
                                                  To_StdLogicVector(INIT_A)  &
                                                  To_StdLogicVector(INIT_9)  &
                                                  To_StdLogicVector(INIT_8)  &
                                                  To_StdLogicVector(INIT_7)  &
                                                  To_StdLogicVector(INIT_6)  &
                                                  To_StdLogicVector(INIT_5)  &
                                                  To_StdLogicVector(INIT_4)  &
                                                  To_StdLogicVector(INIT_3)  &
                                                  To_StdLogicVector(INIT_2)  &
                                                  To_StdLogicVector(INIT_1)  & 
                                                  To_StdLogicVector(INIT_0) ;  

       
  begin

    Violation  := Pviol_WCLK or
                  Tviol_WADDR0_WCLK_posedge or
                  Tviol_WADDR1_WCLK_posedge or
                  Tviol_WADDR2_WCLK_posedge or
                  Tviol_WADDR3_WCLK_posedge or
                  Tviol_WADDR4_WCLK_posedge or
                  Tviol_WADDR5_WCLK_posedge or
                  Tviol_WADDR6_WCLK_posedge or
                  Tviol_WADDR7_WCLK_posedge or
                  Tviol_WADDR8_WCLK_posedge or
                  Tviol_WADDR9_WCLK_posedge or
                  Tviol_WCLKE_WCLK_posedge or
                  Tviol_WE_WCLK_posedge or
                  Tviol_WDATA0_WCLK_posedge or
                  Tviol_WDATA1_WCLK_posedge or
                  Tviol_WDATA2_WCLK_posedge or
                  Tviol_WDATA3_WCLK_posedge or
                  Tviol_WDATA4_WCLK_posedge or
                  Tviol_WDATA5_WCLK_posedge or
                  Tviol_WDATA6_WCLK_posedge or
                  Tviol_WDATA7_WCLK_posedge or
                  Tviol_WDATA8_WCLK_posedge or
                  Tviol_WDATA9_WCLK_posedge or
                  Tviol_WDATA10_WCLK_posedge or
                  Tviol_WDATA11_WCLK_posedge or
                  Tviol_WDATA12_WCLK_posedge or
                  Tviol_WDATA13_WCLK_posedge or
                  Tviol_WDATA14_WCLK_posedge or
                  Tviol_WDATA15_WCLK_posedge or
                  Tviol_MASK0_WCLK_posedge or
                  Tviol_MASK1_WCLK_posedge or
                  Tviol_MASK2_WCLK_posedge or
                  Tviol_MASK3_WCLK_posedge or
                  Tviol_MASK4_WCLK_posedge or
                  Tviol_MASK5_WCLK_posedge or
                  Tviol_MASK6_WCLK_posedge or
                  Tviol_MASK7_WCLK_posedge or
                  Tviol_MASK8_WCLK_posedge or
                  Tviol_MASK9_WCLK_posedge or
                  Tviol_MASK10_WCLK_posedge or
                  Tviol_MASK11_WCLK_posedge or
                  Tviol_MASK12_WCLK_posedge or
                  Tviol_MASK13_WCLK_posedge or
                  Tviol_MASK14_WCLK_posedge or
                  Tviol_MASK15_WCLK_posedge;
 
-------------------------
--  Functionality Section
-------------------------

    WADDR_in <= conv_integer(WADDR_ipd) ;
  
    if (Violation = '1') then
       MEM <= (others => 'X') ;
    elsif ( WCLK_ipd'event and (WCLK_ipd = '1') and (WCLKE_ipd = '1' or WCLKE_ipd = 'H') and (WE_ipd = '1') ) then
       for i in 0 to 15 loop
         if (MASK_ipd(i) = '0') then           
            MEM_temp(16*WADDR_in + i ) := WDATA_ipd(i) ;
         end if ;
       end loop ;
    end if ; 

    MEM <= MEM_temp ;

------------------------
--  Timing Check Section
------------------------
    if (TimingChecksOn) then
      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR0_WCLK_posedge,
        TimingData     => Tmkr_WADDR0_WCLK_posedge,
        TestSignal     => WADDR_ipd(0),
        TestSignalName => "WADDR(0)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(0),
        SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(0),
        HoldLow        => thold_WADDR_WCLK_posedge_posedge(0),
        HoldHigh       => thold_WADDR_WCLK_negedge_posedge(0),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR1_WCLK_posedge,
        TimingData     => Tmkr_WADDR1_WCLK_posedge,
        TestSignal     => WADDR_ipd(1),
        TestSignalName => "WADDR(1)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(1),
        SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(1),
        HoldLow        => thold_WADDR_WCLK_posedge_posedge(1),
        HoldHigh       => thold_WADDR_WCLK_negedge_posedge(1),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR2_WCLK_posedge,
        TimingData     => Tmkr_WADDR2_WCLK_posedge,
        TestSignal     => WADDR_ipd(2),
        TestSignalName => "WADDR(2)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(2),
        SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(2),
        HoldLow        => thold_WADDR_WCLK_posedge_posedge(2),
        HoldHigh       => thold_WADDR_WCLK_negedge_posedge(2),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR3_WCLK_posedge,
        TimingData     => Tmkr_WADDR3_WCLK_posedge,
        TestSignal     => WADDR_ipd(3),
        TestSignalName => "WADDR(3)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(3),
        SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(3),
        HoldLow        => thold_WADDR_WCLK_posedge_posedge(3),
        HoldHigh       => thold_WADDR_WCLK_negedge_posedge(3),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR4_WCLK_posedge,
        TimingData     => Tmkr_WADDR4_WCLK_posedge,
        TestSignal     => WADDR_ipd(4),
        TestSignalName => "WADDR(4)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(4),
        SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(4),
        HoldLow        => thold_WADDR_WCLK_posedge_posedge(4),
        HoldHigh       => thold_WADDR_WCLK_negedge_posedge(4),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR5_WCLK_posedge,
        TimingData     => Tmkr_WADDR5_WCLK_posedge,
        TestSignal     => WADDR_ipd(5),
        TestSignalName => "WADDR(5)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(5),
        SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(5),
        HoldLow        => thold_WADDR_WCLK_posedge_posedge(5),
        HoldHigh       => thold_WADDR_WCLK_negedge_posedge(5),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR6_WCLK_posedge,
        TimingData     => Tmkr_WADDR6_WCLK_posedge,
        TestSignal     => WADDR_ipd(6),
        TestSignalName => "WADDR(6)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(6),
        SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(6),
        HoldLow        => thold_WADDR_WCLK_posedge_posedge(6),
        HoldHigh       => thold_WADDR_WCLK_negedge_posedge(6),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR7_WCLK_posedge,
        TimingData     => Tmkr_WADDR7_WCLK_posedge,
        TestSignal     => WADDR_ipd(7),
        TestSignalName => "WADDR(7)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(7),
        SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(7),
        HoldLow        => thold_WADDR_WCLK_posedge_posedge(7),
        HoldHigh       => thold_WADDR_WCLK_negedge_posedge(7),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);


      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR8_WCLK_posedge,
        TimingData     => Tmkr_WADDR8_WCLK_posedge,
        TestSignal     => WADDR_ipd(8),
        TestSignalName => "WADDR(8)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(8),
        SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(8),
        HoldLow        => thold_WADDR_WCLK_posedge_posedge(8),
        HoldHigh       => thold_WADDR_WCLK_negedge_posedge(8),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WADDR9_WCLK_posedge,
        TimingData     => Tmkr_WADDR9_WCLK_posedge,
        TestSignal     => WADDR_ipd(9),
        TestSignalName => "WADDR(9)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(9),
        SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(9),
        HoldLow        => thold_WADDR_WCLK_posedge_posedge(9),
        HoldHigh       => thold_WADDR_WCLK_negedge_posedge(9),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WCLKE_WCLK_posedge,
        TimingData     => Tmkr_WCLKE_WCLK_posedge,
        TestSignal     => WCLKE_ipd,
        TestSignalName => "WCLKE",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WCLKE_WCLK_posedge_posedge,
        SetupLow       => tsetup_WCLKE_WCLK_negedge_posedge,
        HoldLow        => thold_WCLKE_WCLK_posedge_posedge,
        HoldHigh       => thold_WCLKE_WCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WE_WCLK_posedge,
        TimingData     => Tmkr_WE_WCLK_posedge,
        TestSignal     => WCLK_ipd,
        TestSignalName => "WCLK",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WE_WCLK_posedge_posedge,
        SetupLow       => tsetup_WE_WCLK_negedge_posedge,
        HoldLow        => thold_WE_WCLK_posedge_posedge,
        HoldHigh       => thold_WE_WCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
       VitalSetupHoldCheck (
        Violation      => Tviol_WDATA0_WCLK_posedge,
        TimingData     => Tmkr_WDATA0_WCLK_posedge,
        TestSignal     => WDATA_ipd(0),
        TestSignalName => "WDATA(0)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(0),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(0),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(0),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(0),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA1_WCLK_posedge,
        TimingData     => Tmkr_WDATA1_WCLK_posedge,
        TestSignal     => WDATA_ipd(1),
        TestSignalName => "WDATA(1)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(1),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(1),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(1),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(1),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA2_WCLK_posedge,
        TimingData     => Tmkr_WDATA2_WCLK_posedge,
        TestSignal     => WDATA_ipd(2),
        TestSignalName => "WDATA(2)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(2),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(2),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(2),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(2),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA3_WCLK_posedge,
        TimingData     => Tmkr_WDATA3_WCLK_posedge,
        TestSignal     => WDATA_ipd(3),
        TestSignalName => "WDATA(3)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(3),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(3),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(3),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(3),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA4_WCLK_posedge,
        TimingData     => Tmkr_WDATA4_WCLK_posedge,
        TestSignal     => WDATA_ipd(4),
        TestSignalName => "WDATA(4)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(4),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(4),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(4),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(4),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA5_WCLK_posedge,
        TimingData     => Tmkr_WDATA5_WCLK_posedge,
        TestSignal     => WDATA_ipd(5),
        TestSignalName => "WDATA(5)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(5),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(5),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(5),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(5),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA6_WCLK_posedge,
        TimingData     => Tmkr_WDATA6_WCLK_posedge,
        TestSignal     => WDATA_ipd(6),
        TestSignalName => "WDATA(6)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(6),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(6),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(6),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(6),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA7_WCLK_posedge,
        TimingData     => Tmkr_WDATA7_WCLK_posedge,
        TestSignal     => WDATA_ipd(7),
        TestSignalName => "WDATA(7)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(7),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(7),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(7),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(7),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

       VitalSetupHoldCheck (
        Violation      => Tviol_WDATA8_WCLK_posedge,
        TimingData     => Tmkr_WDATA8_WCLK_posedge,
        TestSignal     => WDATA_ipd(8),
        TestSignalName => "WDATA(8)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(8),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(8),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(8),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(8),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA9_WCLK_posedge,
        TimingData     => Tmkr_WDATA9_WCLK_posedge,
        TestSignal     => WDATA_ipd(9),
        TestSignalName => "WDATA(9)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(9),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(9),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(9),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(9),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA10_WCLK_posedge,
        TimingData     => Tmkr_WDATA10_WCLK_posedge,
        TestSignal     => WDATA_ipd(10),
        TestSignalName => "WDATA(10)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(10),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(10),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(10),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(10),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA11_WCLK_posedge,
        TimingData     => Tmkr_WDATA11_WCLK_posedge,
        TestSignal     => WDATA_ipd(11),
        TestSignalName => "WDATA(11)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(11),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(11),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(11),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(11),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA12_WCLK_posedge,
        TimingData     => Tmkr_WDATA12_WCLK_posedge,
        TestSignal     => WDATA_ipd(12),
        TestSignalName => "WDATA(12)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(12),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(12),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(12),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(12),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA13_WCLK_posedge,
        TimingData     => Tmkr_WDATA13_WCLK_posedge,
        TestSignal     => WDATA_ipd(13),
        TestSignalName => "WDATA(13)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(13),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(13),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(13),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(13),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA14_WCLK_posedge,
        TimingData     => Tmkr_WDATA14_WCLK_posedge,
        TestSignal     => WDATA_ipd(14),
        TestSignalName => "WDATA(14)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(14),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(14),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(14),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(14),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_WDATA15_WCLK_posedge,
        TimingData     => Tmkr_WDATA15_WCLK_posedge,
        TestSignal     => WDATA_ipd(15),
        TestSignalName => "WDATA(15)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(15),
        SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(15),
        HoldLow        => thold_WDATA_WCLK_posedge_posedge(15),
        HoldHigh       => thold_WDATA_WCLK_negedge_posedge(15),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

       VitalSetupHoldCheck (
        Violation      => Tviol_MASK0_WCLK_posedge,
        TimingData     => Tmkr_MASK0_WCLK_posedge,
        TestSignal     => MASK_ipd(0),
        TestSignalName => "MASK(0)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(0),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(0),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(0),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(0),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK1_WCLK_posedge,
        TimingData     => Tmkr_MASK1_WCLK_posedge,
        TestSignal     => MASK_ipd(1),
        TestSignalName => "MASK(1)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(1),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(1),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(1),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(1),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK2_WCLK_posedge,
        TimingData     => Tmkr_MASK2_WCLK_posedge,
        TestSignal     => MASK_ipd(2),
        TestSignalName => "MASK(2)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(2),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(2),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(2),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(2),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK3_WCLK_posedge,
        TimingData     => Tmkr_MASK3_WCLK_posedge,
        TestSignal     => MASK_ipd(3),
        TestSignalName => "MASK(3)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(3),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(3),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(3),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(3),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK4_WCLK_posedge,
        TimingData     => Tmkr_MASK4_WCLK_posedge,
        TestSignal     => MASK_ipd(4),
        TestSignalName => "MASK(4)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(4),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(4),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(4),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(4),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_MASK5_WCLK_posedge,
        TimingData     => Tmkr_MASK5_WCLK_posedge,
        TestSignal     => MASK_ipd(5),
        TestSignalName => "MASK(5)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(5),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(5),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(5),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(5),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_MASK6_WCLK_posedge,
        TimingData     => Tmkr_MASK6_WCLK_posedge,
        TestSignal     => MASK_ipd(6),
        TestSignalName => "MASK(6)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(6),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(6),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(6),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(6),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_MASK7_WCLK_posedge,
        TimingData     => Tmkr_MASK7_WCLK_posedge,
        TestSignal     => MASK_ipd(7),
        TestSignalName => "MASK(7)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(7),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(7),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(7),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(7),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

       VitalSetupHoldCheck (
        Violation      => Tviol_MASK8_WCLK_posedge,
        TimingData     => Tmkr_MASK8_WCLK_posedge,
        TestSignal     => MASK_ipd(8),
        TestSignalName => "MASK(8)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(8),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(8),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(8),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(8),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK9_WCLK_posedge,
        TimingData     => Tmkr_MASK9_WCLK_posedge,
        TestSignal     => MASK_ipd(9),
        TestSignalName => "MASK(9)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(9),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(9),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(9),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(9),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK10_WCLK_posedge,
        TimingData     => Tmkr_MASK10_WCLK_posedge,
        TestSignal     => MASK_ipd(10),
        TestSignalName => "MASK(10)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(10),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(10),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(10),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(10),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK11_WCLK_posedge,
        TimingData     => Tmkr_MASK11_WCLK_posedge,
        TestSignal     => MASK_ipd(11),
        TestSignalName => "MASK(11)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(11),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(11),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(11),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(11),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);        
        
      VitalSetupHoldCheck (
        Violation      => Tviol_MASK12_WCLK_posedge,
        TimingData     => Tmkr_MASK12_WCLK_posedge,
        TestSignal     => MASK_ipd(12),
        TestSignalName => "MASK(12)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(12),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(12),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(12),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(12),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_MASK13_WCLK_posedge,
        TimingData     => Tmkr_MASK13_WCLK_posedge,
        TestSignal     => MASK_ipd(13),
        TestSignalName => "MASK(13)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(13),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(13),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(13),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(13),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_MASK14_WCLK_posedge,
        TimingData     => Tmkr_MASK14_WCLK_posedge,
        TestSignal     => MASK_ipd(14),
        TestSignalName => "MASK(14)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(14),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(14),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(14),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(14),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);

      VitalSetupHoldCheck (
        Violation      => Tviol_MASK15_WCLK_posedge,
        TimingData     => Tmkr_MASK15_WCLK_posedge,
        TestSignal     => MASK_ipd(15),
        TestSignalName => "MASK(15)",
        TestDelay      => 0 ns,
        RefSignal      => WCLK_ipd,
        RefSignalName  => "WCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(15),
        SetupLow       => tsetup_MASK_WCLK_negedge_posedge(15),
        HoldLow        => thold_MASK_WCLK_posedge_posedge(15),
        HoldHigh       => thold_MASK_WCLK_negedge_posedge(15),
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
   

      VitalPeriodPulseCheck (
        Violation      => Pviol_WCLK,
        PeriodData     => PInfo_WCLK,
        TestSignal     => WCLK_ipd,
        TestSignalName => "WCLK",
        TestDelay      => 0 ns,
        Period         => 0 ns,
        PulseWidthHigh => tpw_WCLK_posedge,
        PulseWidthLow  => tpw_WCLK_negedge,
        CheckEnabled   => true,
        HeaderMsg      => "/SB_RAM16K",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);



    end if ;

  end process VITALWriteBehavior;

end SB_RAM16K_V;

------------------------------------
        --- SB_RAM40_16K 
------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;
use IEEE.VITAL_Timing.all;

entity SB_RAM40_16K is

  generic ( 

           TimingChecksOn : boolean := true;
           Xon            : boolean := false;
           MsgOn          : boolean := false;
           
           tipd_RCLK  : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_RCLKE : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_RE    : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_RADDR : VitalDelayArrayType01(12 downto 0) := (others => (0 ns, 0 ns));
           tipd_WCLK  : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_WCLKE : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_WE    : VitalDelayType01                   := ( 0 ns, 0 ns);
           tipd_WADDR : VitalDelayArrayType01(12 downto 0) := (others => (0 ns, 0 ns));
           tipd_MASK  : VitalDelayArrayType01(15 downto 0) := (others => (0 ns, 0 ns));
           tipd_WDATA : VitalDelayArrayType01(15 downto 0) := (others => (0 ns, 0 ns));
		 		
           tpd_RCLK_RDATA : VitalDelayArrayType01(15 downto 0) := (others => (0 ns, 0 ns));
           tpd_RCLK_RDATA_posedge : VitalDelayArrayType01(15 downto 0) := (others => (0 ns, 0 ns));

           tsetup_RADDR_RCLK_negedge_posedge : VitalDelayArrayType(12 downto 0) := (others => 0 ns);
           tsetup_RADDR_RCLK_posedge_posedge : VitalDelayArrayType(12 downto 0) := (others => 0 ns);
           tsetup_RCLKE_RCLK_negedge_posedge : VitalDelayType                   := 0 ns;
           tsetup_RCLKE_RCLK_posedge_posedge : VitalDelayType                   := 0 ns;
           tsetup_RE_RCLK_negedge_posedge    : VitalDelayType                   := 0 ns;
           tsetup_RE_RCLK_posedge_posedge    : VitalDelayType                   := 0 ns;

           tsetup_WADDR_WCLK_negedge_posedge : VitalDelayArrayType(12 downto 0) := (others => 0 ns);
           tsetup_WADDR_WCLK_posedge_posedge : VitalDelayArrayType(12 downto 0) := (others => 0 ns);
           tsetup_WDATA_WCLK_negedge_posedge : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           tsetup_WDATA_WCLK_posedge_posedge : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           tsetup_WCLKE_WCLK_negedge_posedge : VitalDelayType                   := 0 ns;
           tsetup_WCLKE_WCLK_posedge_posedge : VitalDelayType                   := 0 ns;
           tsetup_WE_WCLK_negedge_posedge    : VitalDelayType                   := 0 ns;
           tsetup_WE_WCLK_posedge_posedge    : VitalDelayType                   := 0 ns;
           tsetup_MASK_WCLK_negedge_posedge  : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           tsetup_MASK_WCLK_posedge_posedge  : VitalDelayArrayType(15 downto 0) := (others => 0 ns);

           thold_RADDR_RCLK_negedge_posedge : VitalDelayArrayType(12 downto 0) := (others => 0 ns);
           thold_RADDR_RCLK_posedge_posedge : VitalDelayArrayType(12 downto 0) := (others => 0 ns);
           thold_RCLKE_RCLK_negedge_posedge : VitalDelayType                   := 0 ns;
           thold_RCLKE_RCLK_posedge_posedge : VitalDelayType                   := 0 ns;
           thold_RE_RCLK_negedge_posedge    : VitalDelayType                   := 0 ns;
           thold_RE_RCLK_posedge_posedge    : VitalDelayType                   := 0 ns;

           thold_WADDR_WCLK_negedge_posedge : VitalDelayArrayType(12 downto 0)  := (others => 0 ns);
           thold_WADDR_WCLK_posedge_posedge : VitalDelayArrayType(12 downto 0)  := (others => 0 ns);
           thold_WDATA_WCLK_negedge_posedge : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           thold_WDATA_WCLK_posedge_posedge : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           thold_WCLKE_WCLK_negedge_posedge : VitalDelayType                   := 0 ns;
           thold_WCLKE_WCLK_posedge_posedge : VitalDelayType                   := 0 ns;
           thold_WE_WCLK_negedge_posedge    : VitalDelayType                   := 0 ns;
           thold_WE_WCLK_posedge_posedge    : VitalDelayType                   := 0 ns;
           thold_MASK_WCLK_negedge_posedge  : VitalDelayArrayType(15 downto 0) := (others => 0 ns);
           thold_MASK_WCLK_posedge_posedge  : VitalDelayArrayType(15 downto 0) := (others => 0 ns);

           tpw_RCLK_negedge : VitalDelayType := 0 ns;
           tpw_RCLK_posedge : VitalDelayType := 0 ns;
           tpw_WCLK_negedge : VitalDelayType := 0 ns;
           tpw_WCLK_posedge : VitalDelayType := 0 ns;

	   WRITE_MODE : integer := 0;  -- Configure Write Port as 1024x16 (0)/ 20148x8 (1)/ 4096x4 (2)/ 8192x2 (3)
           READ_MODE  : integer := 0;  -- Configure Read Port as 1024x16 (0)/ 20148x8 (1)/ 4096x4 (2)/ 8192x2 (3)

           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;

          port( 
                RDATA : out std_logic_vector( 15  downto 0) ;
                RCLK  : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'H';
                RADDR : in  std_logic_vector( 12 downto 0) ;
                WCLK  : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'H';
                WADDR : in  std_logic_vector( 12  downto 0) ;
                MASK  : in  std_logic_vector( 15  downto 0) ;
                WDATA : in  std_logic_vector( 15  downto 0)
               );
  
  attribute VITAL_LEVEL0 of SB_RAM40_16K : entity is TRUE;
 
end SB_RAM40_16K;


architecture SB_RAM40_16K_ARCH of SB_RAM40_16K is

  attribute VITAL_LEVEL0 of SB_RAM40_16K_ARCH  : architecture is TRUE;
  
	 component read_data_decoder 
		generic (
			READ_MODE : integer := 0
		);
		port (
			di	 :  in std_logic_vector (15 downto 0);
			ldo	 :  out std_logic_vector (15 downto 0);
			ai	 :  in std_logic_vector (2 downto 0)
		);
	end component;

	component mask_decoder 
		generic (
			WRITE_MODE : integer := 0 
		);
		port (
			mi	 :  in std_logic_vector (15 downto 0);
			mo	 :  out std_logic_vector (15 downto 0);
			ai	 :  in std_logic_vector (2 downto 0)
		);
	end component;

	component write_data_decoder 
		generic (
			WRITE_MODE  : integer := 0
		);
		port (
			di	 : in std_logic_vector(15 downto 0);
			ldo	 : out std_logic_vector (15 downto 0)
		);
	end component;

	component SB_RAM16K 
		generic (
			INIT_0	   : bit_vector;
			INIT_1	   : bit_vector;
			INIT_2	   : bit_vector;
			INIT_3	   : bit_vector;
			INIT_4	   : bit_vector;
			INIT_5	   : bit_vector;
			INIT_6	   : bit_vector;
			INIT_7	   : bit_vector;
			INIT_8	   : bit_vector;
			INIT_9	   : bit_vector;
			INIT_A	   : bit_vector;
			INIT_B	   : bit_vector;
			INIT_C	   : bit_vector;
			INIT_D	   : bit_vector;
			INIT_E	   : bit_vector;
			INIT_F	   : bit_vector;

			INIT_10	   : bit_vector;
			INIT_11	   : bit_vector;
			INIT_12	   : bit_vector;
			INIT_13	   : bit_vector;
			INIT_14	   : bit_vector;
			INIT_15	   : bit_vector;
			INIT_16	   : bit_vector;
			INIT_17	   : bit_vector;
			INIT_18	   : bit_vector;
			INIT_19	   : bit_vector;
			INIT_1A	   : bit_vector;
			INIT_1B	   : bit_vector;
			INIT_1C	   : bit_vector;
			INIT_1D	   : bit_vector;
			INIT_1E	   : bit_vector;
			INIT_1F	   : bit_vector;

			INIT_20	   : bit_vector;
			INIT_21	   : bit_vector;
			INIT_22	   : bit_vector;
			INIT_23	   : bit_vector;
			INIT_24	   : bit_vector;
			INIT_25	   : bit_vector;
			INIT_26	   : bit_vector;
			INIT_27	   : bit_vector;
			INIT_28	   : bit_vector;
			INIT_29	   : bit_vector;
			INIT_2A	   : bit_vector;
			INIT_2B	   : bit_vector;
			INIT_2C	   : bit_vector;
			INIT_2D	   : bit_vector;
			INIT_2E	   : bit_vector;
			INIT_2F	   : bit_vector;

			INIT_30	   : bit_vector;
			INIT_31	   : bit_vector;
			INIT_32	   : bit_vector;
			INIT_33	   : bit_vector;
			INIT_34	   : bit_vector;
			INIT_35	   : bit_vector;
			INIT_36	   : bit_vector;
			INIT_37	   : bit_vector;
			INIT_38	   : bit_vector;
			INIT_39	   : bit_vector;
			INIT_3A	   : bit_vector;
			INIT_3B	   : bit_vector;
			INIT_3C	   : bit_vector;
			INIT_3D	   : bit_vector;
			INIT_3E	   : bit_vector;
			INIT_3F	   : bit_vector
		);
		port (
			RDATA	   : out std_logic_vector(15 downto 0);
			RCLK	   : in std_logic;
			RCLKE	   : in std_logic;
			RE	   : in std_logic;
			RADDR	   : in std_logic_vector(9 downto 0);
			MASK	   : in std_logic_vector(15 downto 0);
			WDATA	   : in std_logic_vector(15 downto 0);
			WCLK	   : in std_logic;
			WCLKE	   : in std_logic;
			WE	   : in std_logic;
			WADDR	   : in std_logic_vector(9 downto 0)
		);
	end component;


	--- VITAL Signals   
	signal RADDR_ipd : std_logic_vector(12 downto 0)  := (others => 'X');   
	signal RCLK_ipd  : std_logic                    := 'X';
	signal RCLKE_ipd : std_logic                    := 'X';
	signal RE_ipd    : std_logic                    := 'X';

	signal WADDR_ipd : std_logic_vector(12 downto 0)  := (others => 'X');
	signal WCLK_ipd  : std_logic                    := 'X';  
	signal WCLKE_ipd : std_logic                    := 'X';
	signal WE_ipd    : std_logic                    := 'X';
	signal MASK_ipd  : std_logic_vector(15 downto 0) := (others => 'X');
	signal WDATA_ipd : std_logic_vector(15 downto 0) := (others => 'X');

        signal RDATA_zd : std_logic_vector(15 downto 0) := (others => 'X');

	---- Function Signals
	signal RD : std_logic_vector(15 downto 0);
	signal WD : std_logic_vector(15 downto 0);
	signal MASK_RAM : std_logic_vector(15 downto 0);

	signal READ_ADDR_HB : std_logic_vector (2 downto 0);
	signal READ_ADDR_LB : std_logic_vector (9 downto 0);
	signal WRITE_ADDR_LB : std_logic_vector (9 downto 0);
	signal WRITE_ADDR_HB : std_logic_vector (2 downto 0);

	signal READ_ADDR_HB_reg : std_logic_vector (2 downto 0); 
	
begin
	---------------------
	--  Input Wire Delay
	---------------------
	WireDelay : block
	begin
	  RADDR_DELAY : for i in 12 downto 0 generate
	     VitalWireDelay (RADDR_ipd(i), RADDR(i), tipd_RADDR(i));
	  end generate RADDR_DELAY;
	  VitalWireDelay (RCLK_ipd, RCLK, tipd_RCLK);
	  VitalWireDelay (RCLKE_ipd, RCLKE, tipd_RCLKE);
	  VitalWireDelay (RE_ipd, RE, tipd_RE);
	  WADDR_DELAY : for i in 12 downto 0 generate
	     VitalWireDelay (WADDR_ipd(i), WADDR(i), tipd_WADDR(i));
	  end generate WADDR_DELAY;
	  VitalWireDelay (WCLK_ipd, WCLK, tipd_WCLK);
	  VitalWireDelay (WCLKE_ipd, WCLKE, tipd_WCLKE);
	  VitalWireDelay (WE_ipd, WE, tipd_WE);
	  MASK_DELAY : for i in 15 downto 0 generate
	     VitalWireDelay (MASK_ipd(i), MASK(i), tipd_MASK(i));
	  end generate MASK_DELAY;
	  WDATA_DELAY : for i in 15 downto 0 generate
	     VitalWireDelay (WDATA_ipd(i), WDATA(i), tipd_WDATA(i));
	  end generate WDATA_DELAY;
	end block;

	VITALBehavior : block
	begin

	---------------------
	--  Timing Checks
	---------------------
	TimingChecks : process (RADDR_ipd, RCLK_ipd, RCLKE_ipd, RE_ipd, WADDR_ipd, WCLK_ipd, WCLKE_ipd, WE_ipd, MASK_ipd, WDATA_ipd)

	variable Tviol_RADDR0_RCLK_posedge : std_logic := '0';
	variable Tviol_RADDR1_RCLK_posedge : std_logic := '0';
	variable Tviol_RADDR2_RCLK_posedge : std_logic := '0';
	variable Tviol_RADDR3_RCLK_posedge : std_logic := '0';
	variable Tviol_RADDR4_RCLK_posedge : std_logic := '0';
	variable Tviol_RADDR5_RCLK_posedge : std_logic := '0';
	variable Tviol_RADDR6_RCLK_posedge : std_logic := '0';
	variable Tviol_RADDR7_RCLK_posedge : std_logic := '0';
	variable Tviol_RADDR8_RCLK_posedge : std_logic := '0';
	variable Tviol_RADDR9_RCLK_posedge : std_logic := '0';
	variable Tviol_RADDR10_RCLK_posedge : std_logic := '0';
	variable Tviol_RADDR11_RCLK_posedge : std_logic := '0';
	variable Tviol_RADDR12_RCLK_posedge : std_logic := '0';
	variable Tviol_RCLKE_RCLK_posedge  : std_logic := '0';
	variable Tviol_RE_RCLK_posedge     : std_logic := '0';

	variable Tmkr_RADDR0_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_RADDR1_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_RADDR2_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_RADDR3_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_RADDR4_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_RADDR5_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_RADDR6_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_RADDR7_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_RADDR8_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_RADDR9_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_RADDR10_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_RADDR11_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_RADDR12_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_RCLKE_RCLK_posedge  : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_RE_RCLK_posedge     : VitalTimingDataType := VitalTimingDataInit;

	variable PViol_RCLK : std_logic := '0';

	variable PInfo_RCLK : VitalPeriodDataType ;

        variable Tviol_WADDR0_WCLK_posedge : std_logic := '0';
        variable Tviol_WADDR1_WCLK_posedge : std_logic := '0';
        variable Tviol_WADDR2_WCLK_posedge : std_logic := '0';
        variable Tviol_WADDR3_WCLK_posedge : std_logic := '0';
        variable Tviol_WADDR4_WCLK_posedge : std_logic := '0';
        variable Tviol_WADDR5_WCLK_posedge : std_logic := '0';
        variable Tviol_WADDR6_WCLK_posedge : std_logic := '0';
        variable Tviol_WADDR7_WCLK_posedge : std_logic := '0';
        variable Tviol_WADDR8_WCLK_posedge : std_logic := '0';
        variable Tviol_WADDR9_WCLK_posedge : std_logic := '0';
        variable Tviol_WADDR10_WCLK_posedge : std_logic := '0';
        variable Tviol_WADDR11_WCLK_posedge : std_logic := '0';
        variable Tviol_WADDR12_WCLK_posedge : std_logic := '0';
        variable Tviol_WCLKE_WCLK_posedge  : std_logic := '0';
        variable Tviol_WE_WCLK_posedge     : std_logic := '0';
        variable Tviol_WDATA0_WCLK_posedge : std_logic := '0';
        variable Tviol_WDATA1_WCLK_posedge : std_logic := '0';
        variable Tviol_WDATA2_WCLK_posedge : std_logic := '0';
        variable Tviol_WDATA3_WCLK_posedge : std_logic := '0';
        variable Tviol_WDATA4_WCLK_posedge : std_logic := '0';
        variable Tviol_WDATA5_WCLK_posedge : std_logic := '0';
        variable Tviol_WDATA6_WCLK_posedge : std_logic := '0';
        variable Tviol_WDATA7_WCLK_posedge : std_logic := '0';
        variable Tviol_WDATA8_WCLK_posedge : std_logic := '0';
        variable Tviol_WDATA9_WCLK_posedge : std_logic := '0';
        variable Tviol_WDATA10_WCLK_posedge : std_logic := '0';
        variable Tviol_WDATA11_WCLK_posedge : std_logic := '0';
        variable Tviol_WDATA12_WCLK_posedge : std_logic := '0';
        variable Tviol_WDATA13_WCLK_posedge : std_logic := '0';
        variable Tviol_WDATA14_WCLK_posedge : std_logic := '0';
        variable Tviol_WDATA15_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK0_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK1_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK2_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK3_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK4_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK5_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK6_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK7_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK8_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK9_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK10_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK11_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK12_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK13_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK14_WCLK_posedge : std_logic := '0';
        variable Tviol_MASK15_WCLK_posedge : std_logic := '0';


        variable Tmkr_WADDR0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WADDR1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WADDR2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WADDR3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WADDR4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WADDR5_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WADDR6_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WADDR7_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WADDR8_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WADDR9_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WADDR10_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WADDR11_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WADDR12_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WCLKE_WCLK_posedge  : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WE_WCLK_posedge     : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA5_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA6_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA7_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA8_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA9_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA10_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA11_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA12_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA13_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA14_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_WDATA15_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK5_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK6_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK7_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK8_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK9_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK10_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK11_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK12_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK13_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK14_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
        variable Tmkr_MASK15_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;

        variable PViol_WCLK : std_logic := '0';

        variable PInfo_WCLK : VitalPeriodDataType := VitalPeriodDataInit;

	variable Violation     : std_logic  := '0';

	begin

	    if (TimingChecksOn) then
	      VitalSetupHoldCheck (
		Violation      => Tviol_RADDR0_RCLK_posedge,
		TimingData     => Tmkr_RADDR0_RCLK_posedge,
		TestSignal     => RADDR_ipd(0),
		TestSignalName => "RADDR(0)",
		TestDelay      => 0 ns,
		RefSignal      => RCLK_ipd,
		RefSignalName  => "RCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(0),
		SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(0),
		HoldLow        => thold_RADDR_RCLK_posedge_posedge(0),
		HoldHigh       => thold_RADDR_RCLK_negedge_posedge(0),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_RADDR1_RCLK_posedge,
		TimingData     => Tmkr_RADDR1_RCLK_posedge,
		TestSignal     => RADDR_ipd(1),
		TestSignalName => "RADDR(1)",
		TestDelay      => 0 ns,
		RefSignal      => RCLK_ipd,
		RefSignalName  => "RCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(1),
		SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(1),
		HoldLow        => thold_RADDR_RCLK_posedge_posedge(1),
		HoldHigh       => thold_RADDR_RCLK_negedge_posedge(1),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_RADDR2_RCLK_posedge,
		TimingData     => Tmkr_RADDR2_RCLK_posedge,
		TestSignal     => RADDR_ipd(2),
		TestSignalName => "RADDR(2)",
		TestDelay      => 0 ns,
		RefSignal      => RCLK_ipd,
		RefSignalName  => "RCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(2),
		SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(2),
		HoldLow        => thold_RADDR_RCLK_posedge_posedge(2),
		HoldHigh       => thold_RADDR_RCLK_negedge_posedge(2),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_RADDR3_RCLK_posedge,
		TimingData     => Tmkr_RADDR3_RCLK_posedge,
		TestSignal     => RADDR_ipd(3),
		TestSignalName => "RADDR(3)",
		TestDelay      => 0 ns,
		RefSignal      => RCLK_ipd,
		RefSignalName  => "RCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(3),
		SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(3),
		HoldLow        => thold_RADDR_RCLK_posedge_posedge(3),
		HoldHigh       => thold_RADDR_RCLK_negedge_posedge(3),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_RADDR4_RCLK_posedge,
		TimingData     => Tmkr_RADDR4_RCLK_posedge,
		TestSignal     => RADDR_ipd(4),
		TestSignalName => "RADDR(4)",
		TestDelay      => 0 ns,
		RefSignal      => RCLK_ipd,
		RefSignalName  => "RCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(4),
		SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(4),
		HoldLow        => thold_RADDR_RCLK_posedge_posedge(4),
		HoldHigh       => thold_RADDR_RCLK_negedge_posedge(4),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_RADDR5_RCLK_posedge,
		TimingData     => Tmkr_RADDR5_RCLK_posedge,
		TestSignal     => RADDR_ipd(5),
		TestSignalName => "RADDR(5)",
		TestDelay      => 0 ns,
		RefSignal      => RCLK_ipd,
		RefSignalName  => "RCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(5),
		SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(5),
		HoldLow        => thold_RADDR_RCLK_posedge_posedge(5),
		HoldHigh       => thold_RADDR_RCLK_negedge_posedge(5),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_RADDR6_RCLK_posedge,
		TimingData     => Tmkr_RADDR6_RCLK_posedge,
		TestSignal     => RADDR_ipd(6),
		TestSignalName => "RADDR(6)",
		TestDelay      => 0 ns,
		RefSignal      => RCLK_ipd,
		RefSignalName  => "RCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(6),
		SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(6),
		HoldLow        => thold_RADDR_RCLK_posedge_posedge(6),
		HoldHigh       => thold_RADDR_RCLK_negedge_posedge(6),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);


	      VitalSetupHoldCheck (
		Violation      => Tviol_RADDR7_RCLK_posedge,
		TimingData     => Tmkr_RADDR7_RCLK_posedge,
		TestSignal     => RADDR_ipd(7),
		TestSignalName => "RADDR(7)",
		TestDelay      => 0 ns,
		RefSignal      => RCLK_ipd,
		RefSignalName  => "RCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(7),
		SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(7),
		HoldLow        => thold_RADDR_RCLK_posedge_posedge(7),
		HoldHigh       => thold_RADDR_RCLK_negedge_posedge(7),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_RADDR8_RCLK_posedge,
		TimingData     => Tmkr_RADDR8_RCLK_posedge,
		TestSignal     => RADDR_ipd(8),
		TestSignalName => "RADDR(8)",
		TestDelay      => 0 ns,
		RefSignal      => RCLK_ipd,
		RefSignalName  => "RCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(8),
		SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(8),
		HoldLow        => thold_RADDR_RCLK_posedge_posedge(8),
		HoldHigh       => thold_RADDR_RCLK_negedge_posedge(8),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_RADDR9_RCLK_posedge,
		TimingData     => Tmkr_RADDR9_RCLK_posedge,
		TestSignal     => RADDR_ipd(9),
		TestSignalName => "RADDR(9)",
		TestDelay      => 0 ns,
		RefSignal      => RCLK_ipd,
		RefSignalName  => "RCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(9),
		SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(9),
		HoldLow        => thold_RADDR_RCLK_posedge_posedge(9),
		HoldHigh       => thold_RADDR_RCLK_negedge_posedge(9),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_RADDR10_RCLK_posedge,
		TimingData     => Tmkr_RADDR10_RCLK_posedge,
		TestSignal     => RADDR_ipd(10),
		TestSignalName => "RADDR(10)",
		TestDelay      => 0 ns,
		RefSignal      => RCLK_ipd,
		RefSignalName  => "RCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(10),
		SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(10),
		HoldLow        => thold_RADDR_RCLK_posedge_posedge(10),
		HoldHigh       => thold_RADDR_RCLK_negedge_posedge(10),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_RADDR11_RCLK_posedge,
		TimingData     => Tmkr_RADDR11_RCLK_posedge,
		TestSignal     => RADDR_ipd(11),
		TestSignalName => "RADDR(11)",
		TestDelay      => 0 ns,
		RefSignal      => RCLK_ipd,
		RefSignalName  => "RCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(11),
		SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(11),
		HoldLow        => thold_RADDR_RCLK_posedge_posedge(11),
		HoldHigh       => thold_RADDR_RCLK_negedge_posedge(11),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_RADDR12_RCLK_posedge,
		TimingData     => Tmkr_RADDR12_RCLK_posedge,
		TestSignal     => RADDR_ipd(12),
		TestSignalName => "RADDR(12)",
		TestDelay      => 0 ns,
		RefSignal      => RCLK_ipd,
		RefSignalName  => "RCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_RADDR_RCLK_posedge_posedge(12),
		SetupLow       => tsetup_RADDR_RCLK_negedge_posedge(12),
		HoldLow        => thold_RADDR_RCLK_posedge_posedge(12),
		HoldHigh       => thold_RADDR_RCLK_negedge_posedge(12),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_RCLKE_RCLK_posedge,
		TimingData     => Tmkr_RCLKE_RCLK_posedge,
		TestSignal     => RCLKE_ipd,
		TestSignalName => "RCLKE",
		TestDelay      => 0 ns,
		RefSignal      => RCLK_ipd,
		RefSignalName  => "RCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_RCLKE_RCLK_posedge_posedge,
		SetupLow       => tsetup_RCLKE_RCLK_negedge_posedge,
		HoldLow        => thold_RCLKE_RCLK_posedge_posedge,
		HoldHigh       => thold_RCLKE_RCLK_negedge_posedge,
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_RE_RCLK_posedge,
		TimingData     => Tmkr_RE_RCLK_posedge,
		TestSignal     => RCLK_ipd,
		TestSignalName => "RCLK",
		TestDelay      => 0 ns,
		RefSignal      => RCLK_ipd,
		RefSignalName  => "RCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_RE_RCLK_posedge_posedge,
		SetupLow       => tsetup_RE_RCLK_negedge_posedge,
		HoldLow        => thold_RE_RCLK_posedge_posedge,
		HoldHigh       => thold_RE_RCLK_negedge_posedge,
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		       

	      VitalPeriodPulseCheck (
		Violation      => Pviol_RCLK,
		PeriodData     => PInfo_RCLK,
		TestSignal     => RCLK_ipd,
		TestSignalName => "RCLK",
		TestDelay      => 0 ns,
		Period         => 0 ns,
		PulseWidthHigh => tpw_RCLK_posedge,
		PulseWidthLow  => tpw_RCLK_negedge,
		CheckEnabled   => true,
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_WADDR0_WCLK_posedge,
		TimingData     => Tmkr_WADDR0_WCLK_posedge,
		TestSignal     => WADDR_ipd(0),
		TestSignalName => "WADDR(0)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(0),
		SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(0),
		HoldLow        => thold_WADDR_WCLK_posedge_posedge(0),
		HoldHigh       => thold_WADDR_WCLK_negedge_posedge(0),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_WADDR1_WCLK_posedge,
		TimingData     => Tmkr_WADDR1_WCLK_posedge,
		TestSignal     => WADDR_ipd(1),
		TestSignalName => "WADDR(1)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(1),
		SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(1),
		HoldLow        => thold_WADDR_WCLK_posedge_posedge(1),
		HoldHigh       => thold_WADDR_WCLK_negedge_posedge(1),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_WADDR2_WCLK_posedge,
		TimingData     => Tmkr_WADDR2_WCLK_posedge,
		TestSignal     => WADDR_ipd(2),
		TestSignalName => "WADDR(2)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(2),
		SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(2),
		HoldLow        => thold_WADDR_WCLK_posedge_posedge(2),
		HoldHigh       => thold_WADDR_WCLK_negedge_posedge(2),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_WADDR3_WCLK_posedge,
		TimingData     => Tmkr_WADDR3_WCLK_posedge,
		TestSignal     => WADDR_ipd(3),
		TestSignalName => "WADDR(3)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(3),
		SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(3),
		HoldLow        => thold_WADDR_WCLK_posedge_posedge(3),
		HoldHigh       => thold_WADDR_WCLK_negedge_posedge(3),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_WADDR4_WCLK_posedge,
		TimingData     => Tmkr_WADDR4_WCLK_posedge,
		TestSignal     => WADDR_ipd(4),
		TestSignalName => "WADDR(4)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(4),
		SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(4),
		HoldLow        => thold_WADDR_WCLK_posedge_posedge(4),
		HoldHigh       => thold_WADDR_WCLK_negedge_posedge(4),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_WADDR5_WCLK_posedge,
		TimingData     => Tmkr_WADDR5_WCLK_posedge,
		TestSignal     => WADDR_ipd(5),
		TestSignalName => "WADDR(5)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(5),
		SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(5),
		HoldLow        => thold_WADDR_WCLK_posedge_posedge(5),
		HoldHigh       => thold_WADDR_WCLK_negedge_posedge(5),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_WADDR6_WCLK_posedge,
		TimingData     => Tmkr_WADDR6_WCLK_posedge,
		TestSignal     => WADDR_ipd(6),
		TestSignalName => "WADDR(6)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(6),
		SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(6),
		HoldLow        => thold_WADDR_WCLK_posedge_posedge(6),
		HoldHigh       => thold_WADDR_WCLK_negedge_posedge(6),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_WADDR7_WCLK_posedge,
		TimingData     => Tmkr_WADDR7_WCLK_posedge,
		TestSignal     => WADDR_ipd(7),
		TestSignalName => "WADDR(7)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(7),
		SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(7),
		HoldLow        => thold_WADDR_WCLK_posedge_posedge(7),
		HoldHigh       => thold_WADDR_WCLK_negedge_posedge(7),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);


	      VitalSetupHoldCheck (
		Violation      => Tviol_WADDR8_WCLK_posedge,
		TimingData     => Tmkr_WADDR8_WCLK_posedge,
		TestSignal     => WADDR_ipd(8),
		TestSignalName => "WADDR(8)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(8),
		SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(8),
		HoldLow        => thold_WADDR_WCLK_posedge_posedge(8),
		HoldHigh       => thold_WADDR_WCLK_negedge_posedge(8),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);


	      VitalSetupHoldCheck (
		Violation      => Tviol_WADDR9_WCLK_posedge,
		TimingData     => Tmkr_WADDR9_WCLK_posedge,
		TestSignal     => WADDR_ipd(9),
		TestSignalName => "WADDR(9)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(9),
		SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(9),
		HoldLow        => thold_WADDR_WCLK_posedge_posedge(9),
		HoldHigh       => thold_WADDR_WCLK_negedge_posedge(9),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);


	      VitalSetupHoldCheck (
		Violation      => Tviol_WADDR10_WCLK_posedge,
		TimingData     => Tmkr_WADDR10_WCLK_posedge,
		TestSignal     => WADDR_ipd(10),
		TestSignalName => "WADDR(10)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(10),
		SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(10),
		HoldLow        => thold_WADDR_WCLK_posedge_posedge(10),
		HoldHigh       => thold_WADDR_WCLK_negedge_posedge(10),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_WADDR11_WCLK_posedge,
		TimingData     => Tmkr_WADDR11_WCLK_posedge,
		TestSignal     => WADDR_ipd(11),
		TestSignalName => "WADDR(11)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(11),
		SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(11),
		HoldLow        => thold_WADDR_WCLK_posedge_posedge(11),
		HoldHigh       => thold_WADDR_WCLK_negedge_posedge(11),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_WADDR12_WCLK_posedge,
		TimingData     => Tmkr_WADDR12_WCLK_posedge,
		TestSignal     => WADDR_ipd(12),
		TestSignalName => "WADDR(12)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WADDR_WCLK_posedge_posedge(12),
		SetupLow       => tsetup_WADDR_WCLK_negedge_posedge(12),
		HoldLow        => thold_WADDR_WCLK_posedge_posedge(12),
		HoldHigh       => thold_WADDR_WCLK_negedge_posedge(12),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_WCLKE_WCLK_posedge,
		TimingData     => Tmkr_WCLKE_WCLK_posedge,
		TestSignal     => WCLKE_ipd,
		TestSignalName => "WCLKE",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WCLKE_WCLK_posedge_posedge,
		SetupLow       => tsetup_WCLKE_WCLK_negedge_posedge,
		HoldLow        => thold_WCLKE_WCLK_posedge_posedge,
		HoldHigh       => thold_WCLKE_WCLK_negedge_posedge,
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_WE_WCLK_posedge,
		TimingData     => Tmkr_WE_WCLK_posedge,
		TestSignal     => WCLK_ipd,
		TestSignalName => "WCLK",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WE_WCLK_posedge_posedge,
		SetupLow       => tsetup_WE_WCLK_negedge_posedge,
		HoldLow        => thold_WE_WCLK_posedge_posedge,
		HoldHigh       => thold_WE_WCLK_negedge_posedge,
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	       VitalSetupHoldCheck (
		Violation      => Tviol_WDATA0_WCLK_posedge,
		TimingData     => Tmkr_WDATA0_WCLK_posedge,
		TestSignal     => WDATA_ipd(0),
		TestSignalName => "WDATA(0)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(0),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(0),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(0),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(0),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_WDATA1_WCLK_posedge,
		TimingData     => Tmkr_WDATA1_WCLK_posedge,
		TestSignal     => WDATA_ipd(1),
		TestSignalName => "WDATA(1)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(1),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(1),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(1),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(1),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_WDATA2_WCLK_posedge,
		TimingData     => Tmkr_WDATA2_WCLK_posedge,
		TestSignal     => WDATA_ipd(2),
		TestSignalName => "WDATA(2)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(2),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(2),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(2),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(2),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_WDATA3_WCLK_posedge,
		TimingData     => Tmkr_WDATA3_WCLK_posedge,
		TestSignal     => WDATA_ipd(3),
		TestSignalName => "WDATA(3)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(3),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(3),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(3),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(3),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_WDATA4_WCLK_posedge,
		TimingData     => Tmkr_WDATA4_WCLK_posedge,
		TestSignal     => WDATA_ipd(4),
		TestSignalName => "WDATA(4)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(4),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(4),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(4),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(4),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_WDATA5_WCLK_posedge,
		TimingData     => Tmkr_WDATA5_WCLK_posedge,
		TestSignal     => WDATA_ipd(5),
		TestSignalName => "WDATA(5)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(5),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(5),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(5),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(5),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_WDATA6_WCLK_posedge,
		TimingData     => Tmkr_WDATA6_WCLK_posedge,
		TestSignal     => WDATA_ipd(6),
		TestSignalName => "WDATA(6)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(6),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(6),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(6),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(6),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_WDATA7_WCLK_posedge,
		TimingData     => Tmkr_WDATA7_WCLK_posedge,
		TestSignal     => WDATA_ipd(7),
		TestSignalName => "WDATA(7)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(7),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(7),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(7),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(7),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	       VitalSetupHoldCheck (
		Violation      => Tviol_WDATA8_WCLK_posedge,
		TimingData     => Tmkr_WDATA8_WCLK_posedge,
		TestSignal     => WDATA_ipd(8),
		TestSignalName => "WDATA(8)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(8),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(8),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(8),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(8),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_WDATA9_WCLK_posedge,
		TimingData     => Tmkr_WDATA9_WCLK_posedge,
		TestSignal     => WDATA_ipd(9),
		TestSignalName => "WDATA(9)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(9),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(9),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(9),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(9),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_WDATA10_WCLK_posedge,
		TimingData     => Tmkr_WDATA10_WCLK_posedge,
		TestSignal     => WDATA_ipd(10),
		TestSignalName => "WDATA(10)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(10),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(10),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(10),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(10),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_WDATA11_WCLK_posedge,
		TimingData     => Tmkr_WDATA11_WCLK_posedge,
		TestSignal     => WDATA_ipd(11),
		TestSignalName => "WDATA(11)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(11),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(11),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(11),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(11),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_WDATA12_WCLK_posedge,
		TimingData     => Tmkr_WDATA12_WCLK_posedge,
		TestSignal     => WDATA_ipd(12),
		TestSignalName => "WDATA(12)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(12),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(12),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(12),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(12),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_WDATA13_WCLK_posedge,
		TimingData     => Tmkr_WDATA13_WCLK_posedge,
		TestSignal     => WDATA_ipd(13),
		TestSignalName => "WDATA(13)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(13),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(13),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(13),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(13),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_WDATA14_WCLK_posedge,
		TimingData     => Tmkr_WDATA14_WCLK_posedge,
		TestSignal     => WDATA_ipd(14),
		TestSignalName => "WDATA(14)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(14),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(14),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(14),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(14),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_WDATA15_WCLK_posedge,
		TimingData     => Tmkr_WDATA15_WCLK_posedge,
		TestSignal     => WDATA_ipd(15),
		TestSignalName => "WDATA(15)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WDATA_WCLK_posedge_posedge(15),
		SetupLow       => tsetup_WDATA_WCLK_negedge_posedge(15),
		HoldLow        => thold_WDATA_WCLK_posedge_posedge(15),
		HoldHigh       => thold_WDATA_WCLK_negedge_posedge(15),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	       VitalSetupHoldCheck (
		Violation      => Tviol_MASK0_WCLK_posedge,
		TimingData     => Tmkr_MASK0_WCLK_posedge,
		TestSignal     => MASK_ipd(0),
		TestSignalName => "MASK(0)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(0),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(0),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(0),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(0),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_MASK1_WCLK_posedge,
		TimingData     => Tmkr_MASK1_WCLK_posedge,
		TestSignal     => MASK_ipd(1),
		TestSignalName => "MASK(1)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(1),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(1),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(1),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(1),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_MASK2_WCLK_posedge,
		TimingData     => Tmkr_MASK2_WCLK_posedge,
		TestSignal     => MASK_ipd(2),
		TestSignalName => "MASK(2)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(2),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(2),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(2),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(2),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_MASK3_WCLK_posedge,
		TimingData     => Tmkr_MASK3_WCLK_posedge,
		TestSignal     => MASK_ipd(3),
		TestSignalName => "MASK(3)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(3),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(3),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(3),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(3),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_MASK4_WCLK_posedge,
		TimingData     => Tmkr_MASK4_WCLK_posedge,
		TestSignal     => MASK_ipd(4),
		TestSignalName => "MASK(4)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(4),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(4),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(4),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(4),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_MASK5_WCLK_posedge,
		TimingData     => Tmkr_MASK5_WCLK_posedge,
		TestSignal     => MASK_ipd(5),
		TestSignalName => "MASK(5)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(5),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(5),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(5),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(5),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_MASK6_WCLK_posedge,
		TimingData     => Tmkr_MASK6_WCLK_posedge,
		TestSignal     => MASK_ipd(6),
		TestSignalName => "MASK(6)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(6),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(6),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(6),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(6),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_MASK7_WCLK_posedge,
		TimingData     => Tmkr_MASK7_WCLK_posedge,
		TestSignal     => MASK_ipd(7),
		TestSignalName => "MASK(7)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(7),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(7),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(7),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(7),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	       VitalSetupHoldCheck (
		Violation      => Tviol_MASK8_WCLK_posedge,
		TimingData     => Tmkr_MASK8_WCLK_posedge,
		TestSignal     => MASK_ipd(8),
		TestSignalName => "MASK(8)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(8),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(8),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(8),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(8),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_MASK9_WCLK_posedge,
		TimingData     => Tmkr_MASK9_WCLK_posedge,
		TestSignal     => MASK_ipd(9),
		TestSignalName => "MASK(9)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(9),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(9),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(9),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(9),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_MASK10_WCLK_posedge,
		TimingData     => Tmkr_MASK10_WCLK_posedge,
		TestSignal     => MASK_ipd(10),
		TestSignalName => "MASK(10)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(10),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(10),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(10),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(10),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_MASK11_WCLK_posedge,
		TimingData     => Tmkr_MASK11_WCLK_posedge,
		TestSignal     => MASK_ipd(11),
		TestSignalName => "MASK(11)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(11),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(11),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(11),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(11),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);        
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_MASK12_WCLK_posedge,
		TimingData     => Tmkr_MASK12_WCLK_posedge,
		TestSignal     => MASK_ipd(12),
		TestSignalName => "MASK(12)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(12),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(12),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(12),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(12),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_MASK13_WCLK_posedge,
		TimingData     => Tmkr_MASK13_WCLK_posedge,
		TestSignal     => MASK_ipd(13),
		TestSignalName => "MASK(13)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(13),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(13),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(13),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(13),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_MASK14_WCLK_posedge,
		TimingData     => Tmkr_MASK14_WCLK_posedge,
		TestSignal     => MASK_ipd(14),
		TestSignalName => "MASK(14)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(14),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(14),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(14),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(14),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_MASK15_WCLK_posedge,
		TimingData     => Tmkr_MASK15_WCLK_posedge,
		TestSignal     => MASK_ipd(15),
		TestSignalName => "MASK(15)",
		TestDelay      => 0 ns,
		RefSignal      => WCLK_ipd,
		RefSignalName  => "WCLK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASK_WCLK_posedge_posedge(15),
		SetupLow       => tsetup_MASK_WCLK_negedge_posedge(15),
		HoldLow        => thold_MASK_WCLK_posedge_posedge(15),
		HoldHigh       => thold_MASK_WCLK_negedge_posedge(15),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
	   

	      VitalPeriodPulseCheck (
		Violation      => Pviol_WCLK,
		PeriodData     => PInfo_WCLK,
		TestSignal     => WCLK_ipd,
		TestSignalName => "WCLK",
		TestDelay      => 0 ns,
		Period         => 0 ns,
		PulseWidthHigh => tpw_WCLK_posedge,
		PulseWidthLow  => tpw_WCLK_negedge,
		CheckEnabled   => true,
		HeaderMsg      => "/SB_RAM40_16K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	    Violation  := Pviol_RCLK or
			  Tviol_RADDR0_RCLK_posedge or
			  Tviol_RADDR1_RCLK_posedge or
			  Tviol_RADDR2_RCLK_posedge or
			  Tviol_RADDR3_RCLK_posedge or
			  Tviol_RADDR4_RCLK_posedge or
			  Tviol_RADDR5_RCLK_posedge or
			  Tviol_RADDR6_RCLK_posedge or
			  Tviol_RADDR7_RCLK_posedge or
			  Tviol_RADDR8_RCLK_posedge or
			  Tviol_RADDR9_RCLK_posedge or
			  Tviol_RADDR10_RCLK_posedge or
			  Tviol_RADDR11_RCLK_posedge or
			  Tviol_RADDR12_RCLK_posedge or
			  Tviol_RCLKE_RCLK_posedge or
			  Tviol_RE_RCLK_posedge or
    			  Pviol_WCLK or
			  Tviol_WADDR0_WCLK_posedge or
			  Tviol_WADDR1_WCLK_posedge or
			  Tviol_WADDR2_WCLK_posedge or
			  Tviol_WADDR3_WCLK_posedge or
			  Tviol_WADDR4_WCLK_posedge or
			  Tviol_WADDR5_WCLK_posedge or
			  Tviol_WADDR6_WCLK_posedge or
			  Tviol_WADDR7_WCLK_posedge or
			  Tviol_WADDR8_WCLK_posedge or
			  Tviol_WADDR9_WCLK_posedge or
			  Tviol_WADDR10_WCLK_posedge or
			  Tviol_WADDR11_WCLK_posedge or
			  Tviol_WADDR12_WCLK_posedge or
			  Tviol_WCLKE_WCLK_posedge or
			  Tviol_WE_WCLK_posedge or
			  Tviol_WDATA0_WCLK_posedge or
			  Tviol_WDATA1_WCLK_posedge or
			  Tviol_WDATA2_WCLK_posedge or
			  Tviol_WDATA3_WCLK_posedge or
			  Tviol_WDATA4_WCLK_posedge or
			  Tviol_WDATA5_WCLK_posedge or
			  Tviol_WDATA6_WCLK_posedge or
			  Tviol_WDATA7_WCLK_posedge or
			  Tviol_WDATA8_WCLK_posedge or
			  Tviol_WDATA9_WCLK_posedge or
			  Tviol_WDATA10_WCLK_posedge or
			  Tviol_WDATA11_WCLK_posedge or
			  Tviol_WDATA12_WCLK_posedge or
			  Tviol_WDATA13_WCLK_posedge or
			  Tviol_WDATA14_WCLK_posedge or
			  Tviol_WDATA15_WCLK_posedge or
			  Tviol_MASK0_WCLK_posedge or
			  Tviol_MASK1_WCLK_posedge or
			  Tviol_MASK2_WCLK_posedge or
			  Tviol_MASK3_WCLK_posedge or
			  Tviol_MASK4_WCLK_posedge or
			  Tviol_MASK5_WCLK_posedge or
			  Tviol_MASK6_WCLK_posedge or
			  Tviol_MASK7_WCLK_posedge or
			  Tviol_MASK8_WCLK_posedge or
			  Tviol_MASK9_WCLK_posedge or
			  Tviol_MASK10_WCLK_posedge or
			  Tviol_MASK11_WCLK_posedge or
			  Tviol_MASK12_WCLK_posedge or
			  Tviol_MASK13_WCLK_posedge or
			  Tviol_MASK14_WCLK_posedge or
			  Tviol_MASK15_WCLK_posedge;

		assert violation = '0'
			report " Incorrect due to Timing Violations\n"
		severity warning;

	    end if ;
    end process TimingChecks;

------------------------
--  BEHAVIOR SECTION
------------------------

	READ_ADDR_HB <= RADDR_ipd(12) & RADDR_ipd(11) & RADDR_ipd(10);
	WRITE_ADDR_HB <= WADDR_ipd(12) & WADDR_ipd(11) & WADDR_ipd(10);
	READ_ADDR_LB <=  RADDR_ipd(9) & RADDR_ipd(8) &  RADDR_ipd(7) & RADDR_ipd(6) & RADDR_ipd(5)& RADDR_ipd(4) & RADDR_ipd(3) & RADDR_ipd(2) & RADDR_ipd(1) & RADDR_ipd(0);
	WRITE_ADDR_LB <= WADDR_ipd(9) & WADDR_ipd(8) &WADDR_ipd(7) & WADDR_ipd(6) & WADDR_ipd(5)& WADDR_ipd(4) & WADDR_ipd(3) & WADDR_ipd(2) & WADDR_ipd(1) & WADDR_ipd(0);

	LatchAddress:process(RCLK_ipd) 
	begin 
		if(RCLK_ipd'event and RCLK_ipd='1') then 
		READ_ADDR_HB_reg <=READ_ADDR_HB;  
		end if; 
	end process LatchAddress;   

	read_data_decoder_inst  : read_data_decoder 
		generic map (
			READ_MODE => READ_MODE
		)
		port map (
			di	=> RD,
			ai	=> READ_ADDR_HB_reg,
			ldo	=> RDATA_zd
		);

	
	write_data_decoder_inst  : write_data_decoder
		generic map (
			WRITE_MODE => WRITE_MODE
		)
		port map (
			di  => WDATA_ipd,
			ldo  => WD
		);

	mask_data_decoder_inst : mask_decoder
		generic map (
			WRITE_MODE => WRITE_MODE
		)
		port map (
			mi  => MASK_ipd,
			mo  => MASK_RAM,
			ai  => WRITE_ADDR_HB
		);
	ram16k_inst : SB_RAM16K
		generic map (
			INIT_0     => INIT_0,
			INIT_1     => INIT_1,
			INIT_2     => INIT_2,
			INIT_3     => INIT_3,
			INIT_4     => INIT_4,
			INIT_5     => INIT_5,
			INIT_6     => INIT_6,
			INIT_7     => INIT_7,
			INIT_8     => INIT_8,
			INIT_9     => INIT_9,
			INIT_A     => INIT_A,
			INIT_B     => INIT_B,
			INIT_C     => INIT_C,
			INIT_D     => INIT_D,
			INIT_E     => INIT_E,
			INIT_F     => INIT_F,

			INIT_10     => INIT_10,
			INIT_11     => INIT_11,
			INIT_12     => INIT_12,
			INIT_13     => INIT_13,
			INIT_14     => INIT_14,
			INIT_15     => INIT_15,
			INIT_16     => INIT_16,
			INIT_17     => INIT_17,
			INIT_18     => INIT_18,
			INIT_19     => INIT_19,
			INIT_1A     => INIT_1A,
			INIT_1B     => INIT_1B,
			INIT_1C     => INIT_1C,
			INIT_1D     => INIT_1D,
			INIT_1E     => INIT_1E,
			INIT_1F     => INIT_1F,

			INIT_20     => INIT_20,
			INIT_21     => INIT_21,
			INIT_22     => INIT_22,
			INIT_23     => INIT_23,
			INIT_24     => INIT_24,
			INIT_25     => INIT_25,
			INIT_26     => INIT_26,
			INIT_27     => INIT_27,
			INIT_28     => INIT_28,
			INIT_29     => INIT_29,
			INIT_2A     => INIT_2A,
			INIT_2B     => INIT_2B,
			INIT_2C     => INIT_2C,
			INIT_2D     => INIT_2D,
			INIT_2E     => INIT_2E,
			INIT_2F     => INIT_2F,

			INIT_30     => INIT_30,
			INIT_31     => INIT_31,
			INIT_32     => INIT_32,
			INIT_33     => INIT_33,
			INIT_34     => INIT_34,
			INIT_35     => INIT_35,
			INIT_36     => INIT_36,
			INIT_37     => INIT_37,
			INIT_38     => INIT_38,
			INIT_39     => INIT_39,
			INIT_3A     => INIT_3A,
			INIT_3B     => INIT_3B,
			INIT_3C     => INIT_3C,
			INIT_3D     => INIT_3D,
			INIT_3E     => INIT_3E,
			INIT_3F     => INIT_3F
		)
		port map (
			RDATA	=> RD,
			RCLK	=> RCLK_ipd,
			RCLKE	=> RCLKE_ipd,
			RE	=> RE_ipd,
			RADDR	=> READ_ADDR_LB,
			MASK	=> MASK_RAM,
			WDATA	=> WD,       
			WCLK	=> WCLK_ipd,
			WCLKE	=> WCLKE_ipd,
			WE	=> WE_ipd,
			WADDR	=> WRITE_ADDR_LB
		);

------------------------
--  Path Delay Section
------------------------
	PathDelay : process(RDATA_zd)

	variable RDATA_GlitchData0  : VitalGlitchDataType;
	variable RDATA_GlitchData1  : VitalGlitchDataType;
	variable RDATA_GlitchData2  : VitalGlitchDataType;
	variable RDATA_GlitchData3  : VitalGlitchDataType;
	variable RDATA_GlitchData4  : VitalGlitchDataType;
	variable RDATA_GlitchData5  : VitalGlitchDataType;
	variable RDATA_GlitchData6  : VitalGlitchDataType;
	variable RDATA_GlitchData7  : VitalGlitchDataType;
	variable RDATA_GlitchData8  : VitalGlitchDataType;
	variable RDATA_GlitchData9  : VitalGlitchDataType;
	variable RDATA_GlitchData10 : VitalGlitchDataType;
	variable RDATA_GlitchData11 : VitalGlitchDataType;
	variable RDATA_GlitchData12 : VitalGlitchDataType;
	variable RDATA_GlitchData13 : VitalGlitchDataType;
	variable RDATA_GlitchData14 : VitalGlitchDataType;
	variable RDATA_GlitchData15 : VitalGlitchDataType;
	begin
	    VitalPathDelay01 (
	      OutSignal     => RDATA(0),
	      GlitchData    => RDATA_GlitchData0,
	      OutSignalName => "RDATA(0)",
	      OutTemp       => RDATA_zd(0),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(0), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => RDATA(1),
	      GlitchData    => RDATA_GlitchData1,
	      OutSignalName => "RDATA(1)",
	      OutTemp       => RDATA_zd(1),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(1), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => RDATA(2),
	      GlitchData    => RDATA_GlitchData2,
	      OutSignalName => "RDATA(2)",
	      OutTemp       => RDATA_zd(2),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(2), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => RDATA(3),
	      GlitchData    => RDATA_GlitchData3,
	      OutSignalName => "RDATA(3)",
	      OutTemp       => RDATA_zd(3),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(3), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => RDATA(4),
	      GlitchData    => RDATA_GlitchData4,
	      OutSignalName => "RDATA(4)",
	      OutTemp       => RDATA_zd(4),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(4), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => RDATA(5),
	      GlitchData    => RDATA_GlitchData5,
	      OutSignalName => "RDATA(5)",
	      OutTemp       => RDATA_zd(5),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(5), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => RDATA(6),
	      GlitchData    => RDATA_GlitchData6,
	      OutSignalName => "RDATA(6)",
	      OutTemp       => RDATA_zd(6),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(6), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => RDATA(7),
	      GlitchData    => RDATA_GlitchData7,
	      OutSignalName => "RDATA(7)",
	      OutTemp       => RDATA_zd(7),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(7), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => RDATA(8),
	      GlitchData    => RDATA_GlitchData8,
	      OutSignalName => "RDATA(8)",
	      OutTemp       => RDATA_zd(8),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(8), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => RDATA(9),
	      GlitchData    => RDATA_GlitchData9,
	      OutSignalName => "RDATA(9)",
	      OutTemp       => RDATA_zd(9),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(9), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => RDATA(10),
	      GlitchData    => RDATA_GlitchData10,
	      OutSignalName => "RDATA(10)",
	      OutTemp       => RDATA_zd(10),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(10), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => RDATA(11),
	      GlitchData    => RDATA_GlitchData11,
	      OutSignalName => "RDATA(11)",
	      OutTemp       => RDATA_zd(11),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(11), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => RDATA(12),
	      GlitchData    => RDATA_GlitchData12,
	      OutSignalName => "RDATA(12)",
	      OutTemp       => RDATA_zd(12),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(12), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => RDATA(13),
	      GlitchData    => RDATA_GlitchData13,
	      OutSignalName => "RDATA(13)",
	      OutTemp       => RDATA_zd(13),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(13), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => RDATA(14),
	      GlitchData    => RDATA_GlitchData14,
	      OutSignalName => "RDATA(14)",
	      OutTemp       => RDATA_zd(14),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(14), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => RDATA(15),
	      GlitchData    => RDATA_GlitchData15,
	      OutSignalName => "RDATA(15)",
	      OutTemp       => RDATA_zd(15),
	      Paths         => (0 => (RCLK_ipd'last_event, tpd_RCLK_RDATA(15), true)),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	end process;

	end block;

end SB_RAM40_16K_ARCH;   --- SB_RAM40_16K


---------------------------------------
	--- SB_RAM40_16KNR
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM40_16KNR is

  generic ( 
	   WRITE_MODE : integer := 0; -- Configure Write Port as 1024x16 (0)/ 20148x8 (1)/ 4096x4 (2)/ 8192x2 (3) 
  	   READ_MODE  : integer := 0;  -- Configure Read Port as 1024x16 (0)/ 20148x8 (1)/ 4096x4 (2)/ 8192x2 (3)

           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 15  downto 0) ;
                RCLKN : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'H';
                RADDR : in  std_logic_vector( 12  downto 0) ;
                WCLK  : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'H';
                WADDR : in  std_logic_vector( 12  downto 0) ;
                MASK  : in  std_logic_vector( 15  downto 0) ;
                WDATA : in  std_logic_vector( 15  downto 0)
               );
  
end SB_RAM40_16KNR;

architecture SB_RAM40_16KNR_ARCH of SB_RAM40_16KNR is

	component SB_RAM40_16K
		generic (
			WRITE_MODE : integer;
			READ_MODE  : integer;
			INIT_0	   : bit_vector;
			INIT_1	   : bit_vector;
			INIT_2	   : bit_vector;
			INIT_3	   : bit_vector;
			INIT_4	   : bit_vector;
			INIT_5	   : bit_vector;
			INIT_6	   : bit_vector;
			INIT_7	   : bit_vector;
			INIT_8	   : bit_vector;
			INIT_9	   : bit_vector;
			INIT_A	   : bit_vector;
			INIT_B	   : bit_vector;
			INIT_C	   : bit_vector;
			INIT_D	   : bit_vector;
			INIT_E	   : bit_vector;
			INIT_F	   : bit_vector;

			INIT_10	   : bit_vector;
			INIT_11	   : bit_vector;
			INIT_12	   : bit_vector;
			INIT_13	   : bit_vector;
			INIT_14	   : bit_vector;
			INIT_15	   : bit_vector;
			INIT_16	   : bit_vector;
			INIT_17	   : bit_vector;
			INIT_18	   : bit_vector;
			INIT_19	   : bit_vector;
			INIT_1A	   : bit_vector;
			INIT_1B	   : bit_vector;
			INIT_1C	   : bit_vector;
			INIT_1D	   : bit_vector;
			INIT_1E	   : bit_vector;
			INIT_1F	   : bit_vector;

			INIT_20	   : bit_vector;
			INIT_21	   : bit_vector;
			INIT_22	   : bit_vector;
			INIT_23	   : bit_vector;
			INIT_24	   : bit_vector;
			INIT_25	   : bit_vector;
			INIT_26	   : bit_vector;
			INIT_27	   : bit_vector;
			INIT_28	   : bit_vector;
			INIT_29   : bit_vector;
			INIT_2A	   : bit_vector;
			INIT_2B	   : bit_vector;
			INIT_2C	   : bit_vector;
			INIT_2D	   : bit_vector;
			INIT_2E	   : bit_vector;
			INIT_2F	   : bit_vector;
			
			INIT_30	   : bit_vector;
			INIT_31	   : bit_vector;
			INIT_32	   : bit_vector;
			INIT_33	   : bit_vector;
			INIT_34	   : bit_vector;
			INIT_35	   : bit_vector;
			INIT_36	   : bit_vector;
			INIT_37	   : bit_vector;
			INIT_38	   : bit_vector;
			INIT_39	   : bit_vector;
			INIT_3A	   : bit_vector;
			INIT_3B	   : bit_vector;
			INIT_3C	   : bit_vector;
			INIT_3D	   : bit_vector;
			INIT_3E	   : bit_vector;
			INIT_3F	   : bit_vector
		);
		port (
			RDATA	   : out std_logic_vector(15 downto 0);
			RCLK	   : in std_logic;
			RCLKE	   : in std_logic;
			RE	   : in std_logic;
			RADDR	   : in std_logic_vector(12 downto 0);
			MASK	   : in std_logic_vector(15 downto 0);
			WDATA	   : in std_logic_vector(15 downto 0);
			WCLK	   : in std_logic;
			WCLKE	   : in std_logic;
			WE	   : in std_logic;
			WADDR	   : in std_logic_vector(12 downto 0)
		);
	end component;

	signal RCLK : std_logic;

begin
	RCLK <= not(RCLKN);
	ram40mh_16k_nr_inst : SB_RAM40_16K
		generic map (
			WRITE_MODE => WRITE_MODE,
			READ_MODE  => READ_MODE,
			INIT_0     => INIT_0,
			INIT_1     => INIT_1,
			INIT_2     => INIT_2,
			INIT_3     => INIT_3,
			INIT_4     => INIT_4,
			INIT_5     => INIT_5,
			INIT_6     => INIT_6,
			INIT_7     => INIT_7,
			INIT_8     => INIT_8,
			INIT_9     => INIT_9,
			INIT_A     => INIT_A,
			INIT_B     => INIT_B,
			INIT_C     => INIT_C,
			INIT_D     => INIT_D,
			INIT_E     => INIT_E,
			INIT_F     => INIT_F,

			INIT_10     => INIT_10,
			INIT_11     => INIT_11,
			INIT_12     => INIT_12,
			INIT_13     => INIT_13,
			INIT_14     => INIT_14,
			INIT_15     => INIT_15,
			INIT_16     => INIT_16,
			INIT_17     => INIT_17,
			INIT_18     => INIT_18,
			INIT_19     => INIT_19,
			INIT_1A     => INIT_1A,
			INIT_1B     => INIT_1B,
			INIT_1C     => INIT_1C,
			INIT_1D     => INIT_1D,
			INIT_1E     => INIT_1E,
			INIT_1F     => INIT_1F,

			INIT_20     => INIT_20,
			INIT_21     => INIT_21,
			INIT_22     => INIT_22,
			INIT_23     => INIT_23,
			INIT_24     => INIT_24,
			INIT_25     => INIT_25,
			INIT_26     => INIT_26,
			INIT_27     => INIT_27,
			INIT_28     => INIT_28,
			INIT_29     => INIT_29,
			INIT_2A     => INIT_2A,
			INIT_2B     => INIT_2B,
			INIT_2C     => INIT_2C,
			INIT_2D     => INIT_2D,
			INIT_2E     => INIT_2E,
			INIT_2F     => INIT_2F,

			INIT_30     => INIT_30,
			INIT_31     => INIT_31,
			INIT_32     => INIT_32,
			INIT_33     => INIT_33,
			INIT_34     => INIT_34,
			INIT_35     => INIT_35,
			INIT_36     => INIT_36,
			INIT_37     => INIT_37,
			INIT_38     => INIT_38,
			INIT_39     => INIT_39,
			INIT_3A     => INIT_3A,
			INIT_3B     => INIT_3B,
			INIT_3C     => INIT_3C,
			INIT_3D     => INIT_3D,
			INIT_3E     => INIT_3E,
			INIT_3F     => INIT_3F
		)
		port map (
			RDATA	=> RDATA,
			RCLK	=> RCLK,
			RCLKE	=> RCLKE,
			RE	=> RE,
			RADDR	=> RADDR,
			MASK	=> MASK,
			WDATA	=> WDATA,
			WCLK	=> WCLK,
			WCLKE	=> WCLKE,
			WE	=> WE,
			WADDR	=> WADDR
		);

end SB_RAM40_16KNR_ARCH;   --- SB_RAM40_16KNR


---------------------------------------
	--- SB_RAM40_16KNW
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM40_16KNW is

  generic ( 
	   WRITE_MODE : integer := 0; -- Configure Write Port as 1024x16 (0)/ 20148x8 (1)/ 4096x4 (2)/ 8192x2 (3) 
	   READ_MODE  : integer := 0;  -- Configure Read Port as 1024x16 (0)/ 20148x8 (1)/ 4096x4 (2)/ 8192x2 (3)

           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 15  downto 0) ;
                RCLK  : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'H';
                RADDR : in  std_logic_vector( 12  downto 0) ;
                WCLKN : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'H';
                WADDR : in  std_logic_vector( 12  downto 0) ;
                MASK  : in  std_logic_vector( 15  downto 0) ;
                WDATA : in  std_logic_vector( 15  downto 0)
               );
  
  
end SB_RAM40_16KNW;

architecture SB_RAM40_16KNW_ARCH of SB_RAM40_16KNW is
	
	component SB_RAM40_16K
		generic (
			WRITE_MODE : integer;
			READ_MODE  : integer;
			INIT_0	   : bit_vector;
			INIT_1	   : bit_vector;
			INIT_2	   : bit_vector;
			INIT_3	   : bit_vector;
			INIT_4	   : bit_vector;
			INIT_5	   : bit_vector;
			INIT_6	   : bit_vector;
			INIT_7	   : bit_vector;
			INIT_8	   : bit_vector;
			INIT_9	   : bit_vector;
			INIT_A	   : bit_vector;
			INIT_B	   : bit_vector;
			INIT_C	   : bit_vector;
			INIT_D	   : bit_vector;
			INIT_E	   : bit_vector;
			INIT_F	   : bit_vector;

			INIT_10	   : bit_vector;
			INIT_11	   : bit_vector;
			INIT_12	   : bit_vector;
			INIT_13	   : bit_vector;
			INIT_14	   : bit_vector;
			INIT_15	   : bit_vector;
			INIT_16	   : bit_vector;
			INIT_17	   : bit_vector;
			INIT_18	   : bit_vector;
			INIT_19	   : bit_vector;
			INIT_1A	   : bit_vector;
			INIT_1B	   : bit_vector;
			INIT_1C	   : bit_vector;
			INIT_1D	   : bit_vector;
			INIT_1E	   : bit_vector;
			INIT_1F	   : bit_vector;

			INIT_20	   : bit_vector;
			INIT_21	   : bit_vector;
			INIT_22	   : bit_vector;
			INIT_23	   : bit_vector;
			INIT_24	   : bit_vector;
			INIT_25	   : bit_vector;
			INIT_26	   : bit_vector;
			INIT_27	   : bit_vector;
			INIT_28	   : bit_vector;
			INIT_29   : bit_vector;
			INIT_2A	   : bit_vector;
			INIT_2B	   : bit_vector;
			INIT_2C	   : bit_vector;
			INIT_2D	   : bit_vector;
			INIT_2E	   : bit_vector;
			INIT_2F	   : bit_vector;
			
			INIT_30	   : bit_vector;
			INIT_31	   : bit_vector;
			INIT_32	   : bit_vector;
			INIT_33	   : bit_vector;
			INIT_34	   : bit_vector;
			INIT_35	   : bit_vector;
			INIT_36	   : bit_vector;
			INIT_37	   : bit_vector;
			INIT_38	   : bit_vector;
			INIT_39	   : bit_vector;
			INIT_3A	   : bit_vector;
			INIT_3B	   : bit_vector;
			INIT_3C	   : bit_vector;
			INIT_3D	   : bit_vector;
			INIT_3E	   : bit_vector;
			INIT_3F	   : bit_vector
		);
		port (
			RDATA	   : out std_logic_vector(15 downto 0);
			RCLK	   : in std_logic;
			RCLKE	   : in std_logic;
			RE	   : in std_logic;
			RADDR	   : in std_logic_vector(12 downto 0);
			MASK	   : in std_logic_vector(15 downto 0);
			WDATA	   : in std_logic_vector(15 downto 0);
			WCLK	   : in std_logic;
			WCLKE	   : in std_logic;
			WE	   : in std_logic;
			WADDR	   : in std_logic_vector(12 downto 0)
		);
	end component;

	signal WCLK : std_logic;

begin
	WCLK <= not(WCLKN);
	ram40mh_16k_nw_inst : SB_RAM40_16K
		generic map (
			WRITE_MODE => WRITE_MODE,
			READ_MODE  => READ_MODE,
			INIT_0     => INIT_0,
			INIT_1     => INIT_1,
			INIT_2     => INIT_2,
			INIT_3     => INIT_3,
			INIT_4     => INIT_4,
			INIT_5     => INIT_5,
			INIT_6     => INIT_6,
			INIT_7     => INIT_7,
			INIT_8     => INIT_8,
			INIT_9     => INIT_9,
			INIT_A     => INIT_A,
			INIT_B     => INIT_B,
			INIT_C     => INIT_C,
			INIT_D     => INIT_D,
			INIT_E     => INIT_E,
			INIT_F     => INIT_F,

			INIT_10     => INIT_10,
			INIT_11     => INIT_11,
			INIT_12     => INIT_12,
			INIT_13     => INIT_13,
			INIT_14     => INIT_14,
			INIT_15     => INIT_15,
			INIT_16     => INIT_16,
			INIT_17     => INIT_17,
			INIT_18     => INIT_18,
			INIT_19     => INIT_19,
			INIT_1A     => INIT_1A,
			INIT_1B     => INIT_1B,
			INIT_1C     => INIT_1C,
			INIT_1D     => INIT_1D,
			INIT_1E     => INIT_1E,
			INIT_1F     => INIT_1F,

			INIT_20     => INIT_20,
			INIT_21     => INIT_21,
			INIT_22     => INIT_22,
			INIT_23     => INIT_23,
			INIT_24     => INIT_24,
			INIT_25     => INIT_25,
			INIT_26     => INIT_26,
			INIT_27     => INIT_27,
			INIT_28     => INIT_28,
			INIT_29     => INIT_29,
			INIT_2A     => INIT_2A,
			INIT_2B     => INIT_2B,
			INIT_2C     => INIT_2C,
			INIT_2D     => INIT_2D,
			INIT_2E     => INIT_2E,
			INIT_2F     => INIT_2F,

			INIT_30     => INIT_30,
			INIT_31     => INIT_31,
			INIT_32     => INIT_32,
			INIT_33     => INIT_33,
			INIT_34     => INIT_34,
			INIT_35     => INIT_35,
			INIT_36     => INIT_36,
			INIT_37     => INIT_37,
			INIT_38     => INIT_38,
			INIT_39     => INIT_39,
			INIT_3A     => INIT_3A,
			INIT_3B     => INIT_3B,
			INIT_3C     => INIT_3C,
			INIT_3D     => INIT_3D,
			INIT_3E     => INIT_3E,
			INIT_3F     => INIT_3F
		)
		port map (
			RDATA	=> RDATA,
			RCLK	=> RCLK,
			RCLKE	=> RCLKE,
			RE	=> RE,
			RADDR	=> RADDR,
			MASK	=> MASK,
			WDATA	=> WDATA,
			WCLK	=> WCLK,
			WCLKE	=> WCLKE,
			WE	=> WE,
			WADDR	=> WADDR
		);
end SB_RAM40_16KNW_ARCH;   --- SB_RAM40_16KNW



---------------------------------------
	--- SB_RAM40_16KNRNW
---------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
USE IEEE.numeric_std.ALL;

entity SB_RAM40_16KNRNW is

  generic ( 
	   WRITE_MODE : integer := 0; -- Configure Write Port as 1024x16 (0)/ 20148x8 (1)/ 4096x4 (2)/ 8192x2 (3) 
           READ_MODE  : integer := 0;  -- Configure Read Port as 1024x16 (0)/ 20148x8 (1)/ 4096x4 (2)/ 8192x2 (3)

           INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"; 

           INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
           INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000" 
            ) ;
          port( 
                RDATA : out std_logic_vector( 15  downto 0) ;
                RCLKN : in  std_logic ;
                RCLKE : in  std_logic := 'H';
                RE    : in  std_logic := 'H';
                RADDR : in  std_logic_vector( 12  downto 0) ;
                WCLKN : in  std_logic ;
                WCLKE : in  std_logic := 'H';
                WE    : in  std_logic := 'H';
                WADDR : in  std_logic_vector( 12  downto 0) ;
                MASK  : in  std_logic_vector( 15  downto 0) ;
                WDATA : in  std_logic_vector( 15  downto 0)
               );
  
  
end SB_RAM40_16KNRNW;

architecture SB_RAM40_16KNRNW_ARCH of SB_RAM40_16KNRNW is

	component SB_RAM40_16K
		generic (
			WRITE_MODE : integer;
			READ_MODE  : integer;
			INIT_0	   : bit_vector;
			INIT_1	   : bit_vector;
			INIT_2	   : bit_vector;
			INIT_3	   : bit_vector;
			INIT_4	   : bit_vector;
			INIT_5	   : bit_vector;
			INIT_6	   : bit_vector;
			INIT_7	   : bit_vector;
			INIT_8	   : bit_vector;
			INIT_9	   : bit_vector;
			INIT_A	   : bit_vector;
			INIT_B	   : bit_vector;
			INIT_C	   : bit_vector;
			INIT_D	   : bit_vector;
			INIT_E	   : bit_vector;
			INIT_F	   : bit_vector;

			INIT_10	   : bit_vector;
			INIT_11	   : bit_vector;
			INIT_12	   : bit_vector;
			INIT_13	   : bit_vector;
			INIT_14	   : bit_vector;
			INIT_15	   : bit_vector;
			INIT_16	   : bit_vector;
			INIT_17	   : bit_vector;
			INIT_18	   : bit_vector;
			INIT_19	   : bit_vector;
			INIT_1A	   : bit_vector;
			INIT_1B	   : bit_vector;
			INIT_1C	   : bit_vector;
			INIT_1D	   : bit_vector;
			INIT_1E	   : bit_vector;
			INIT_1F	   : bit_vector;

			INIT_20	   : bit_vector;
			INIT_21	   : bit_vector;
			INIT_22	   : bit_vector;
			INIT_23	   : bit_vector;
			INIT_24	   : bit_vector;
			INIT_25	   : bit_vector;
			INIT_26	   : bit_vector;
			INIT_27	   : bit_vector;
			INIT_28	   : bit_vector;
			INIT_29   : bit_vector;
			INIT_2A	   : bit_vector;
			INIT_2B	   : bit_vector;
			INIT_2C	   : bit_vector;
			INIT_2D	   : bit_vector;
			INIT_2E	   : bit_vector;
			INIT_2F	   : bit_vector;
			
			INIT_30	   : bit_vector;
			INIT_31	   : bit_vector;
			INIT_32	   : bit_vector;
			INIT_33	   : bit_vector;
			INIT_34	   : bit_vector;
			INIT_35	   : bit_vector;
			INIT_36	   : bit_vector;
			INIT_37	   : bit_vector;
			INIT_38	   : bit_vector;
			INIT_39	   : bit_vector;
			INIT_3A	   : bit_vector;
			INIT_3B	   : bit_vector;
			INIT_3C	   : bit_vector;
			INIT_3D	   : bit_vector;
			INIT_3E	   : bit_vector;
			INIT_3F	   : bit_vector
		);
		port (
			RDATA	   : out std_logic_vector(15 downto 0);
			RCLK	   : in std_logic;
			RCLKE	   : in std_logic;
			RE	   : in std_logic;
			RADDR	   : in std_logic_vector(12 downto 0);
			MASK	   : in std_logic_vector(15 downto 0);
			WDATA	   : in std_logic_vector(15 downto 0);
			WCLK	   : in std_logic;
			WCLKE	   : in std_logic;
			WE	   : in std_logic;
			WADDR	   : in std_logic_vector(12 downto 0)
		);
	end component;

	signal RCLK : std_logic; 
	signal WCLK : std_logic;

begin
	RCLK <= not(RCLKN); 
	WCLK <= not(WCLKN);
	ram40mh_16k_nrnw_inst : SB_RAM40_16K
		generic map (
			WRITE_MODE => WRITE_MODE,
			READ_MODE  => READ_MODE,
			INIT_0     => INIT_0,
			INIT_1     => INIT_1,
			INIT_2     => INIT_2,
			INIT_3     => INIT_3,
			INIT_4     => INIT_4,
			INIT_5     => INIT_5,
			INIT_6     => INIT_6,
			INIT_7     => INIT_7,
			INIT_8     => INIT_8,
			INIT_9     => INIT_9,
			INIT_A     => INIT_A,
			INIT_B     => INIT_B,
			INIT_C     => INIT_C,
			INIT_D     => INIT_D,
			INIT_E     => INIT_E,
			INIT_F     => INIT_F,

			INIT_10     => INIT_10,
			INIT_11     => INIT_11,
			INIT_12     => INIT_12,
			INIT_13     => INIT_13,
			INIT_14     => INIT_14,
			INIT_15     => INIT_15,
			INIT_16     => INIT_16,
			INIT_17     => INIT_17,
			INIT_18     => INIT_18,
			INIT_19     => INIT_19,
			INIT_1A     => INIT_1A,
			INIT_1B     => INIT_1B,
			INIT_1C     => INIT_1C,
			INIT_1D     => INIT_1D,
			INIT_1E     => INIT_1E,
			INIT_1F     => INIT_1F,

			INIT_20     => INIT_20,
			INIT_21     => INIT_21,
			INIT_22     => INIT_22,
			INIT_23     => INIT_23,
			INIT_24     => INIT_24,
			INIT_25     => INIT_25,
			INIT_26     => INIT_26,
			INIT_27     => INIT_27,
			INIT_28     => INIT_28,
			INIT_29     => INIT_29,
			INIT_2A     => INIT_2A,
			INIT_2B     => INIT_2B,
			INIT_2C     => INIT_2C,
			INIT_2D     => INIT_2D,
			INIT_2E     => INIT_2E,
			INIT_2F     => INIT_2F,

			INIT_30     => INIT_30,
			INIT_31     => INIT_31,
			INIT_32     => INIT_32,
			INIT_33     => INIT_33,
			INIT_34     => INIT_34,
			INIT_35     => INIT_35,
			INIT_36     => INIT_36,
			INIT_37     => INIT_37,
			INIT_38     => INIT_38,
			INIT_39     => INIT_39,
			INIT_3A     => INIT_3A,
			INIT_3B     => INIT_3B,
			INIT_3C     => INIT_3C,
			INIT_3D     => INIT_3D,
			INIT_3E     => INIT_3E,
			INIT_3F     => INIT_3F
		)
		port map (
			RDATA	=> RDATA,
			RCLK	=> RCLK,
			RCLKE	=> RCLKE,
			RE	=> RE,
			RADDR	=> RADDR,
			MASK	=> MASK,
			WDATA	=> WDATA,
			WCLK	=> WCLK,
			WCLKE	=> WCLKE,
			WE	=> WE,
			WADDR	=> WADDR
		);

end SB_RAM40_16KNRNW_ARCH;   --- SB_RAM40_16KNRNW

-----------------------------------------------------
	--- END iCE40MH RAM  Primitives
-----------------------------------------------------


----------------------------------------------------------------------------
--					preio_physical
----------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity	preio_physical	is

	port	(
			bs_en		:	in	std_logic;		--JTAG enable           
			shift		:	in	std_logic;		--JTAG shift            
			tclk		:	in	std_logic;		--JTAG clock            
			update		:	in	std_logic;		--JTAG update           
			sdi			:	in	std_logic;		--JTAG serial data in   
			mode		:	in	std_logic;		--JTAG mode             
			hiz_b		:	in	std_logic;		--JTAG high X control   
			sdo			:	out	std_logic;		--JTAG serial data out  
			dout1		:	out	std_logic;		--Normal Input cell output 1
			dout0		:	out	std_logic;		--Normal Input cell output 0
			ddr1		:	in	std_logic;		--Normal Output cell input 1
			ddr0		:	in	std_logic;		--Normal Output cell input 0
			oepin		:	in	std_logic;		--Normal Ouput-Enable       
			hold		:	in	std_logic;		--Normal Input cell control 
			rstio		:	in	std_logic;		--Normal Input cell reset   
			inclk		:	in	std_logic;		--Normal Input cell clock   
			outclk		:	in	std_logic;		--Normal Output cell clock  
			cbit		:	in	std_logic_vector (5 downto 0);	--Configurion bits   
			padin		:	in	std_logic;		--PAD input          
			padout		:	out	std_logic;		--PAD output         
			padoen		:	out	std_logic 		--PAD output enable  
			);

end preio_physical;

	
architecture preio_physical_v of preio_physical is
--  attribute VITAL_LEVEL0 of
  --  preio_physical_v : architecture is true;
	
	signal	padin_n1,inclk_n2,padin_n3	:	std_logic;
	signal	in_MUX_n4	:	std_logic;
	signal	hold_AND2	:	std_logic;
	signal	ddr0_n11	:	std_logic;
	signal	outclk_n12	:	std_logic;
	signal	ddr1_n13	:	std_logic;
	signal	n14			:	std_logic;
	signal	dout_reg_0_n	:	std_logic;
	signal	Reg_or_Wire_N17	:	std_logic;
	signal	n18			:	std_logic;
	signal	n19			:	std_logic;
	signal	tristate	:	std_logic;
	signal	outclk_n22	:	std_logic;
	signal	n26			:	std_logic;
	signal	oen_n_n24	:	std_logic;
	signal	jtag_update_n30	:	std_logic;
	signal	din_reg_0	:	std_logic;
	signal  din_reg_1	:	std_logic;
	signal	dout_reg_0	:	std_logic;
	signal	dout_reg_1	:	std_logic;
	signal	tristate_q	:	std_logic;
	signal	jtag_oe_reg	:	std_logic;
	signal	temp1,temp2		:	std_logic_vector (1 downto 0);
	signal	dout_0		:	std_logic;		--	wire for port signal usage
begin
	jtag_update_n30	<=	not	(bs_en and (not update));
	
	sdo		<=	din_reg_0;
	dout1 	<= 	din_reg_1;
--------------------------------------------------------------	
	padin_n1_i	:	process	(dout_reg_0, padin, shift)
				begin
					if	(shift='1')	then
						padin_n1	<=	dout_reg_0;
					else
						padin_n1	<=	padin;
					end if;
				end	process;
	
	inclk_n2_i	:	process	(bs_en, tclk, inclk)
				begin
					if	(bs_en='1')	then
						inclk_n2	<=	tclk;
					else
						inclk_n2	<=	inclk;
					end if;
				end process;

	din_reg_0_i	:	process	(inclk_n2, rstio)
				begin
					if	(rstio='1')	then
						din_reg_0	<=	'0';
					elsif	(inclk_n2 'event and inclk_n2='1') then
						din_reg_0	<=	padin_n1;
					end if;
				end process;
-------------------------------------------------------------				
	padin_n3_i	:	process	(bs_en, din_reg_0, padin)
				begin
					if	(bs_en='1')	then
						padin_n3	<=	din_reg_0;
					else
						padin_n3	<=	padin;
					end if;
				end	process;
	
	din_reg_1_i	:	process	(inclk_n2, rstio)
				begin
					if	(rstio='1')	then
						din_reg_1	<=	'0';
					elsif	(inclk_n2 'event and inclk_n2='0') then
						if	(jtag_update_n30='1')	then
							din_reg_1	<=	padin_n3;
						end if;
					end if;
				end process;
--------------------------------------------------------------	
	hold_AND2 <= cbit(1) and hold;

   	--Input MUX   	
	temp1	<=	hold_AND2 & cbit(0);

	in_MUX_n4_i	:	process	(temp1, dout_0, din_reg_0, padin)
   				begin
   					case	temp1 is
   					when	"00"	=>
   						in_MUX_n4 <= din_reg_0;
   					when	"01"	=>
   						in_MUX_n4 <= padin;
   					when	"10"	=>
   						in_MUX_n4 <= dout_0;
   					when	"11"	=>
   						in_MUX_n4 <= dout_0;
   					when others 	=>
   						in_MUX_n4 <= '0';
   					end case;
   				end process;

------------------------dout0 generate------------------------------
	dout_0_i	:	process	(mode, din_reg_1, in_MUX_n4)
			begin
				if	(mode='1')	then
					dout_0	<=	din_reg_1;
				else
					dout_0	<=	in_MUX_n4;
				end if;
			end process;
	
	dout0	<=	dout_0;
--------------------------------------------------------------------	
	--Output Register
	
	dout_reg_0_i	:	process	(outclk_n12, rstio)
				begin
					if	(rstio='1')	then
						dout_reg_0	<=	'0';
					elsif	(outclk_n12 'event and outclk_n12='1') then
						dout_reg_0	<=	ddr0_n11;
					end if;
				end process;

	--Muxes for Output registers
	
	dout_reg_0_n 	<= not dout_reg_0;
	n19 			<= not (outclk_n12 or cbit(2));
	
	Reg_or_Wire_N17_i	:	process	(cbit(2), dout_reg_0_n, ddr0)
					begin
						if	(cbit(2)='1')	then
							Reg_or_Wire_N17	<=	dout_reg_0_n;
						else
							Reg_or_Wire_N17	<=	ddr0;
						end if;
					end process;
	
	n18_i				:	process	(n19, dout_reg_1, dout_reg_0)
					begin
						if	(n19='1')	then
							n18	<=	dout_reg_1;
						else
							n18	<=	dout_reg_0;
						end if;
					end process;

	n14_i				:	process	(cbit(3), Reg_or_Wire_N17, n18)	
					begin
						if	(cbit(3)='1')	then
							n14	<=	Reg_or_Wire_N17;
						else
							n14	<=	n18;
						end if;
					end process;
					
	padout_i			:	process	(mode, dout_reg_1, n14)
					begin
						if	(mode='1')	then
							padout	<=	dout_reg_1;
						else
							padout	<=	n14;
						end if;
					end process;

	--JTAG Assigns
	
	ddr0_n11_i		:	process	(shift, tristate_q, ddr0)
					begin
						if	(shift='1')	then
							ddr0_n11	<=	tristate_q;
						else
							ddr0_n11	<=	ddr0;
						end if;
					end process;

	outclk_n12_i		:	process	(bs_en, tclk, outclk)
					begin
						if	(bs_en='1')	then
							outclk_n12	<=	tclk;
						else
							outclk_n12	<=	outclk;
						end if;
					end process;
					
	ddr1_n13_i		:	process	(bs_en, dout_reg_0, ddr1)
					begin
						if	(bs_en='1')	then
							ddr1_n13	<=	dout_reg_0;
						else
							ddr1_n13	<=	ddr1;
						end if;
					end process;

	--JTAG register 
	dout_reg_1_i		:	process	(outclk_n12, rstio)
					begin
						if	(rstio='1')	then
							dout_reg_1	<=	'0';
						elsif	(outclk_n12 'event and outclk_n12='0') then
							dout_reg_1	<=	ddr1_n13;
						end if;
					end process;
					
----------------------------------------------------------------------------
--
--	Output Enable Logic
--
-----------------------------------------------------------------------------
	--OE Tristate Register
	tristate_i	:	process	(shift, sdi, oepin)
				begin
					if	(shift='1')	then
						tristate	<=	sdi;
					else
						tristate	<=	oepin;
					end if;
				end process;

	tristate_q_i	:	process	(outclk_n22, rstio)
				begin
					if	(rstio='1')	then
						tristate_q	<=	'0';
					elsif	(outclk_n22 'event and outclk_n22 = '1') then
						tristate_q	<=	tristate;
					end if;
				end process;
				
	--JTAG register
	outclk_n22_i	:	process	(bs_en, tclk, outclk)
				begin
					if	(bs_en='1')	then
						outclk_n22	<=	tclk;
					else
						outclk_n22	<=	outclk;
					end if;
				end process;
	
	jtag_oe_reg_i	:	process	(outclk_n22, rstio)
				begin
					if	(rstio='1')	then
						jtag_oe_reg	<=	'0';
					elsif	(outclk_n22 'event and outclk_n22 ='0') then
						if	(jtag_update_n30='1')	then
							jtag_oe_reg	<=	padin_n3;
						end if;
					end if;
				end process;
	
   	temp2	<=	cbit(5) & cbit(4); 
  	--	oen_n_n24_i	:	process	(cbit(5),cbit(4), oepin, tristate_q) 
  	oen_n_n24_i	:	process	(temp2, oepin, tristate_q) 
  					begin 
  						--case	cbit(5) & cbit(4) is 
  						case	temp2 is 
  							when	"00"	=> 
  							oen_n_n24	<=	'0'; 
  							when	"01"	=> 
  							oen_n_n24	<=	'1'; 
  							when	"10"	=> 
  							oen_n_n24	<=	oepin; 
  							when	"11"	=>
   							oen_n_n24	<=	tristate_q; 
   							when others		=> 
   							oen_n_n24	<=	'0'; 
   						end case; 
   					end process;
	
	n26_i			:	process	(mode, jtag_oe_reg, oen_n_n24)
				begin
					if	(mode='1')	then
						n26	<=	jtag_oe_reg;
					else
						n26	<=	oen_n_n24;
					end if;
				end process;

	padoen <= not (hiz_b and n26);
	
end preio_physical_v;



------------------------------------------------------------------------
--					SB_IO
------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
--library	work;
use	work.std_logic_SBT.all;

entity	SB_IO is

	generic (
			NEG_TRIGGER : bit						:=	'0';
			PIN_TYPE	: bit_vector (5 downto 0)	:=	"000000";
			PULLUP		: bit						:=	'0';
			IO_STANDARD	: string					:=	"SB_LVCMOS"
			);
	port 
		(
		D_OUT_1 		    : in std_logic;
		D_OUT_0 		    : in std_logic;
		CLOCK_ENABLE		: in std_logic;
		LATCH_INPUT_VALUE	: in std_logic;
		INPUT_CLK			: in std_logic;
		
		D_IN_1				: out std_logic;
		D_IN_0				: out std_logic;
		OUTPUT_ENABLE		: in std_logic	:='H';
		OUTPUT_CLK			: in std_logic;
		PACKAGE_PIN			: inout	std_ulogic
		); 
		
end SB_IO ;

architecture SB_IO_V of SB_IO is

	component	preio_physical
	port	(
			hold	:	in 	std_logic;
			rstio	:	in	std_logic;
			bs_en	:	in	std_logic;
			shift	:	in	std_logic;
			tclk	:	in	std_logic;
			inclk	:	in	std_logic;
			outclk	:	in	std_logic;
			update	:	in	std_logic;
			oepin	:	in	std_logic;
			sdi		:	in	std_logic;
			mode	:	in	std_logic;
			hiz_b	:	in	std_logic;
			sdo		:	out	std_logic;
			dout1	:	out	std_logic;
			dout0	:	out	std_logic;
			ddr1	:	in	std_logic;
			ddr0	:	in	std_logic;
			padin	:	in	std_logic;
			padout	:	out	std_logic;
			padoen	:	out	std_logic;
			cbit	:	in	std_logic_vector	(5 downto 0)
			);
	end component;

	signal	inclk_n, outclk_n, inclk, outclk,sdo	:	std_logic;
	
	signal	bs_en	:	std_logic	:='0';	--Boundary scan enable           
	signal	shift	:	std_logic	:='0';	--Boundary scan shift            
	signal	tclk	:	std_logic	:='0';	--Boundary scan clock            
	signal	update	:	std_logic	:='0';	--Boundary scan update           
	signal	sdi		:	std_logic	:='0';	--Boundary scan serial data in   
	signal	mode	:	std_logic	:='0';	--Boundary scan mode             
	signal	hiz_b	:	std_logic	:='1';	--Boundary scan Tristate control 
	
	signal	pin_cbit:	std_logic_vector(5 downto 0);
	signal	neg_trig:	std_logic;
	signal	pull_up	:	std_logic;
	signal	hold,oepin,padoen,padout,padin	:	std_logic;
	signal INCLKE_sync , OUTCLKE_sync  	: std_logic;
begin
	
	pin_cbit	<=	TO_STDLOGICVECTOR	(PIN_TYPE);
	neg_trig	<=	TO_STDLOGIC	(NEG_TRIGGER);
	pull_up		<=	TO_STDLOGIC	(PULLUP);

	inclk_n	<= 	INPUT_CLK xor neg_trig;
	outclk_n<=	OUTPUT_CLK xor neg_trig;
--	inclk	<=	inclk_n and CLOCK_ENABLE;
--	outclk	<=	outclk_n and CLOCK_ENABLE;

	process(inclk_n , CLOCK_ENABLE) is
         begin
                if(inclk_n ='0') then
                        INCLKE_sync  <= CLOCK_ENABLE;
                else
                        INCLKE_sync <= INCLKE_sync;
                end if ;
        end process;

        process(outclk_n , CLOCK_ENABLE) is
        begin
                if(outclk_n ='0') then
                        OUTCLKE_sync  <= CLOCK_ENABLE;
                else
                        OUTCLKE_sync <= OUTCLKE_sync;
                end if ;
        end process;

        inclk <= (inclk_n and INCLKE_sync);
        outclk <= (outclk_n and OUTCLKE_sync);
	
	hold	<=	LATCH_INPUT_VALUE;
	oepin	<=	OUTPUT_ENABLE;
	
	PACKAGE_PIN_i	:	process	(padoen, padout, PACKAGE_PIN)
	begin
		padin	<=	PACKAGE_PIN;
		if	(padoen='1') then
			PACKAGE_PIN	<=	'Z';
		else
			PACKAGE_PIN	<=	padout;
		end if;
	end process;
-----------------------------------------------------------------	
	preio_physical_i	:	preio_physical
	port map	(
				hold	=>	hold,
				rstio	=>	'0',
				bs_en	=>	bs_en,
				shift	=>	shift,
				tclk	=>	tclk,
				inclk	=>	inclk,
				outclk	=>	outclk,
				update	=>	update,
				oepin	=>	oepin,
				sdi		=>	sdi,
				mode	=>	mode,
				hiz_b	=>	hiz_b,
				sdo		=>	sdo,
				dout1	=>	D_IN_1,
				dout0	=>	D_IN_0,
				ddr1	=>	D_OUT_1,
				ddr0	=>	D_OUT_0,
				padin	=>	padin,
				padout	=>	padout,
				padoen	=>	padoen,
				cbit	=>	pin_cbit
				);
end	SB_IO_V;

----------------------------------------------------------------------
--					SB_GB_IO
----------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
--library	work;
use	work.std_logic_SBT.all;

entity	SB_GB_IO is
	generic	(
			NEG_TRIGGER : bit						:=	'0';
			PIN_TYPE	: bit_vector (5 downto 0)	:=	"000000";
			PULLUP		: bit						:=	'0';
			IO_STANDARD	: string					:=	"SB_LVCMOS"
			);
			
	port	(
			PACKAGE_PIN			:	inout	std_ulogic;
			LATCH_INPUT_VALUE	:	in		std_logic;
			CLOCK_ENABLE        :	in		std_logic;
			INPUT_CLK           :	in		std_logic;
			OUTPUT_CLK          :	in		std_logic;
			OUTPUT_ENABLE		: in std_logic	:='H';
			D_OUT_1             :	in		std_logic;
			D_OUT_0             :	in		std_logic;
			D_IN_1              :	out		std_logic;
			D_IN_0              :	out		std_logic;
			GLOBAL_BUFFER_OUTPUT:	out		std_logic
			);
end SB_GB_IO;

architecture SB_GB_IO_V of SB_GB_IO is

	component	preio_physical
	port	(
			hold	:	in 	std_logic;
			rstio	:	in	std_logic;
			bs_en	:	in	std_logic;
			shift	:	in	std_logic;
			tclk	:	in	std_logic;
			inclk	:	in	std_logic;
			outclk	:	in	std_logic;
			update	:	in	std_logic;
			oepin	:	in	std_logic;
			sdi		:	in	std_logic;
			mode	:	in	std_logic;
			hiz_b	:	in	std_logic;
			sdo		:	out	std_logic;
			dout1	:	out	std_logic;
			dout0	:	out	std_logic;
			ddr1	:	in	std_logic;
			ddr0	:	in	std_logic;
			padin	:	in	std_logic;
			padout	:	out	std_logic;
			padoen	:	out	std_logic;
			cbit	:	in	std_logic_vector	(5 downto 0)
			);
	end component;
	
	signal	inclk_n,outclk_n,inclk,outclk,sdo	:	std_logic;
	
	signal	bs_en	:	std_logic	:='0';	--Boundary scan enable           
	signal	shift	:	std_logic	:='0';	--Boundary scan shift            
	signal	tclk	:	std_logic	:='0';	--Boundary scan clock            
	signal	update	:	std_logic	:='0';	--Boundary scan update           
	signal	sdi		:	std_logic	:='0';	--Boundary scan serial data in   
	signal	mode	:	std_logic	:='0';	--Boundary scan mode             
	signal	hiz_b	:	std_logic	:='1';	--Boundary scan Tristate control 
	
	signal	hold,oepin,padoen,padout,padin	:	std_logic;
	
	signal	neg_trig:	std_logic;
	signal	pull_up	:	std_logic;
	signal	pin_cbit:	std_logic_vector(5 downto 0);
	signal INCLKE_sync, OUTCLKE_sync : std_logic; 
	
begin
	
	neg_trig	<=	TO_STDLOGIC	(NEG_TRIGGER);
	pin_cbit	<=	TO_STDLOGICVECTOR	(PIN_TYPE);
	pull_up		<=	TO_STDLOGIC	(PULLUP);

	inclk_n	<= 	INPUT_CLK xor neg_trig;
	outclk_n	<=	OUTPUT_CLK xor neg_trig;
--	inclk	<=	inclk_n and CLOCK_ENABLE;
--	outclk	<=	outclk_n and CLOCK_ENABLE;

	process(inclk_n , CLOCK_ENABLE) is
         begin
                if(inclk_n ='0') then
                        INCLKE_sync  <= CLOCK_ENABLE;
                else
                        INCLKE_sync <= INCLKE_sync;
                end if ;
        end process;

        process(outclk_n , CLOCK_ENABLE) is
        begin
                if(outclk_n ='0') then
                        OUTCLKE_sync  <= CLOCK_ENABLE;
                else
                        OUTCLKE_sync <= OUTCLKE_sync;
                end if ;
        end process;

        inclk <= (inclk_n and INCLKE_sync);
        outclk <= (outclk_n and OUTCLKE_sync);
	
	hold	<=	LATCH_INPUT_VALUE;
	oepin	<=	OUTPUT_ENABLE;
	
	PACKAGE_PIN_i	:	process	(padoen, padout, PACKAGE_PIN)
	begin
		padin	<=	PACKAGE_PIN;
		if	(padoen='1') then
			PACKAGE_PIN	<=	'Z';
		else
			PACKAGE_PIN	<=	padout;
		end if;
	end process;
	
	GLOBAL_BUFFER_OUTPUT	<=	padin;
-----------------------------------------------------------------	

	preio_physical_i	:	preio_physical
	port map	(
				hold	=>	hold,
				rstio	=>	'0',
				bs_en	=>	bs_en,
				shift	=>	shift,
				tclk	=>	tclk,
				inclk	=>	inclk,
				outclk	=>	outclk,
				update	=>	update,
				oepin	=>	oepin,
				sdi		=>	sdi,
				mode	=>	mode,
				hiz_b	=>	hiz_b,
				sdo		=>	sdo,
				dout1	=>	D_IN_1,
				dout0	=>	D_IN_0,
				ddr1	=>	D_OUT_1,
				ddr0	=>	D_OUT_0,
				padin	=>	padin,
				padout	=>	padout,
				padoen	=>	padoen,
				cbit	=>	pin_cbit
				);
end	SB_GB_IO_V;

-----------------------------------------------------------------
--					SB_GB
-----------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
--library	work;
use	work.std_logic_SBT.all;

entity	SB_GB	is

port	(
		GLOBAL_BUFFER_OUTPUT			:	out	std_logic;
		USER_SIGNAL_TO_GLOBAL_BUFFER	:	in	std_logic
		);

end	SB_GB;

architecture	SB_GB_V of SB_GB is
begin
	GLOBAL_BUFFER_OUTPUT	<=	USER_SIGNAL_TO_GLOBAL_BUFFER;
end SB_GB_V;




library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity	SB_WARMBOOT	is
port	(
		BOOT	:	in	std_logic;
		S1		:	in	std_logic;
		S0		:	in	std_logic
		);

end SB_WARMBOOT;

-----------------------------------------------------------
--				SB_IO_DS
------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
--library	work;
use	work.std_logic_SBT.all;

	--Differential signaling IO
entity	SB_IO_DS	is
	generic	(
			NEG_TRIGGER : bit						:=	'0';
			PIN_TYPE	: bit_vector (5 downto 0)	:=	"000000";
			IO_STANDARD	: string					:=	"SB_LVDS_OUTPUT"
			);

	port	(
			D_OUT_1			:	in	std_logic;	-- Input output 1 
			D_OUT_0			:	in	std_logic;	-- Input output 0 
			CLOCK_ENABLE	:	in	std_logic;	-- Clock enables NEW - common to in/out clocks 
			D_IN_1			:	out	std_logic;	-- Output input 1
			D_IN_0			:	out	std_logic;	-- Output input 0
			OUTPUT_ENABLE		: in std_logic	:='H';	-- Ouput-Enable 
			LATCH_INPUT_VALUE	:	in	std_logic;	-- Input control 
			INPUT_CLK		:	in	std_logic;	-- Input clock 
			OUTPUT_CLK		:	in	std_logic;  -- Output clock
			PACKAGE_PIN		:	inout	std_ulogic;	-- User's package pin - 'PAD' output  
			PACKAGE_PIN_B	:	inout	std_ulogic	-- User's package pin - 'PAD' output  
			);

end SB_IO_DS;

architecture SB_IO_DS_V of SB_IO_DS is
	--	signals
---------------------
	signal	inclk_n,outclk_n,inclk,outclk,sdo	:	std_logic;
	
	signal	bs_en	:	std_logic	:='0';	--Boundary scan enable           
	signal	shift	:	std_logic	:='0';	--Boundary scan shift            
	signal	tclk	:	std_logic	:='0';	--Boundary scan clock            
	signal	update	:	std_logic	:='0';	--Boundary scan update           
	signal	sdi		:	std_logic	:='0';	--Boundary scan serial data in   
	signal	mode	:	std_logic	:='0';	--Boundary scan mode             
	signal	hiz_b	:	std_logic	:='1';	--Boundary scan Tristate control 
	
	signal	hold,oepin	:	std_logic;	--The required package pin type must be set when io_macro is instantiated.
	signal	padoen, padout, padin	:	std_logic;
	
	signal	pin_cbit:	std_logic_vector(5 downto 0);
	signal	neg_trig:	std_logic;
	
	--	component preio_physical
	component	preio_physical
	port	(
			hold	:	in 	std_logic;
			rstio	:	in	std_logic;
			bs_en	:	in	std_logic;
			shift	:	in	std_logic;
			tclk	:	in	std_logic;
			inclk	:	in	std_logic;
			outclk	:	in	std_logic;
			update	:	in	std_logic;
			oepin	:	in	std_logic;
			sdi		:	in	std_logic;
			mode	:	in	std_logic;
			hiz_b	:	in	std_logic;
			sdo		:	out	std_logic;
			dout1	:	out	std_logic;
			dout0	:	out	std_logic;
			ddr1	:	in	std_logic;
			ddr0	:	in	std_logic;
			padin	:	in	std_logic;
			padout	:	out	std_logic;
			padoen	:	out	std_logic;
			cbit	:	in	std_logic_vector	(5 downto 0)
			);
	end component;

	signal INCLKE_sync,OUTCLKE_sync : std_logic; 
begin
	neg_trig	<=	TO_STDLOGIC	(NEG_TRIGGER);
	pin_cbit	<=	TO_STDLOGICVECTOR	(PIN_TYPE);
	

	inclk_n	<= 	INPUT_CLK xor neg_trig;
	outclk_n	<=	OUTPUT_CLK xor neg_trig;
--	inclk	<=	inclk_n and CLOCK_ENABLE;
--	outclk	<=	outclk_n and CLOCK_ENABLE;

	process(inclk_n , CLOCK_ENABLE) is
         begin
                if(inclk_n ='0') then
                        INCLKE_sync  <= CLOCK_ENABLE;
                else
                        INCLKE_sync <= INCLKE_sync;
                end if ;
        end process;

        process(outclk_n , CLOCK_ENABLE) is
        begin
                if(outclk_n ='0') then
                        OUTCLKE_sync  <= CLOCK_ENABLE;
                else
                        OUTCLKE_sync <= OUTCLKE_sync;
                end if ;
        end process;

        inclk <= (inclk_n and INCLKE_sync);
        outclk <= (outclk_n and OUTCLKE_sync);	
	hold	<=	LATCH_INPUT_VALUE;
	oepin	<=	OUTPUT_ENABLE;
	
	PACKAGE_PIN_i	:	process	(padoen, padout)
	begin
		if	(padoen='1') then
			PACKAGE_PIN	<=	'Z';
		else
			PACKAGE_PIN	<=	padout;
		end if;
	end process;
	
	padin <= PACKAGE_PIN ;
	
	PACKAGE_PIN_B_i	:	process	(padoen, padout)
	begin
		if	(padoen='1') then
			PACKAGE_PIN_B	<=	'Z';
		else
			PACKAGE_PIN_B	<=	not padout;
		end if;
	end process;

	hold	<= LATCH_INPUT_VALUE;
	oepin 	<= OUTPUT_ENABLE;

--	preio_physical_i
	preio_physical_i	:	preio_physical
	port map	(
				hold	=>	hold,
				rstio	=>	'0',
				bs_en	=>	bs_en,
				shift	=>	shift,
				tclk	=>	tclk,
				inclk	=>	inclk,
				outclk	=>	outclk,
				update	=>	update,
				oepin	=>	oepin,
				sdi		=>	sdi,
				mode	=>	mode,
				hiz_b	=>	hiz_b,
				sdo		=>	sdo,
				dout1	=>	D_IN_1,
				dout0	=>	D_IN_0,
				ddr1	=>	D_OUT_1,
				ddr0	=>	D_OUT_0,
				padin	=>	padin,
				padout	=>	padout,
				padoen	=>	padoen,
				cbit	=>	pin_cbit
				);

end SB_IO_DS_V; 

------------------------------------------------------------------------
--					SB_IO
------------------------------------------------------------------------
--
--library ieee;
--use ieee.std_logic_1164.all;
--use ieee.std_logic_arith.all;
--use ieee.std_logic_unsigned.all;
--use IEEE.Vital_Primitives.all;
--use IEEE.VITAL_Timing.all;
----library	work;
--use	work.std_logic_SBT.all;
--
--
--
--entity	SB_IO is
--
--	generic (
--			NEG_TRIGGER : bit						:=	'0';
--			PIN_TYPE	: bit_vector (5 downto 0)	:=	"010000";
--			PULLUP		: bit						:=	'0';
--			IO_STANDARD	: string					:=	"SB_LVCMOS";
--			----------------------------------------------------------------------------------
--			--VITAL PARAMETER
--			---------------------------------------------------------------------------------
--			TimingChecksOn  : boolean := true;
--			Xon   : boolean := true;
--            MsgOn : boolean := false;
--			--- VITAL path delay
--			tipd_D_OUT_1       : VitalDelayType01 := (0 ns, 0 ns);
--            tipd_D_OUT_0       : VitalDelayType01 := (0 ns, 0 ns);
--            tipd_CLOCK_ENABLE        : VitalDelayType01 := (0 ns, 0 ns);
--            tipd_LATCH_INPUT_VALUE       : VitalDelayType01 := (0 ns, 0 ns);
--            tipd_INPUT_CLK        : VitalDelayType01 := (0 ns, 0 ns);
--			tipd_OUTPUT_ENABLE       : VitalDelayType01 := (0 ns, 0 ns);
--            tipd_OUTPUT_CLK       : VitalDelayType01 := (0 ns, 0 ns);
--			tipd_PACKAGE_PIN      : VitalDelayType01 := (0 ns, 0 ns);
--            --- VITAL path delay
--            tpd_PACKAGE_PIN_D_IN_0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
--            tpd_PACKAGE_PIN_D_IN_1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
--            tpd_D_OUT_0_PACKAGE_PIN : VitalDelayType01 := (0.000 ns, 0.000 ns);
--			tpd_D_OUT_1_PACKAGE_PIN : VitalDelayType01 := (0.000 ns, 0.000 ns);
--            tpd_OUTPUT_ENABLE_PACKAGE_PIN : VitalDelayType01 := (0.000 ns, 0.000 ns);
--            tpd_LATCH_INPUT_VALUE_D_IN_0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
--			tpd_LATCH_INPUT_VALUE_D_IN_1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
--			--  VITAL clk-to-output path delay
--			tpd_INPUT_CLK_D_IN_0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
--            tpd_INPUT_CLK_D_IN_1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
--			tpd_OUTPUT_CLK_PACKAGE_PIN : VitalDelayType01 := (0.000 ns, 0.000 ns);
--			--- VITAL setup time
--			tsetup_CLOCK_ENABLE_INPUT_CLK_negedge_posedge    : VitalDelayType                   := 0 ns;
--            tsetup_CLOCK_ENABLE_INPUT_CLK_posedge_posedge    : VitalDelayType                   := 0 ns;
--            tsetup_PACKAGE_PIN_INPUT_CLK_negedge_posedge : VitalDelayType                   := 0 ns;
--            tsetup_PACKAGE_PIN_INPUT_CLK_posedge_posedge : VitalDelayType                   := 0 ns;
--            tsetup_PACKAGE_PIN_INPUT_CLK_posedge_negedge : VitalDelayType                   := 0 ns;
--            tsetup_PACKAGE_PIN_INPUT_CLK_negedge_negedge : VitalDelayType                   := 0 ns;
--            tsetup_CLOCK_ENABLE_OUTPUT_CLK_negedge_posedge   : VitalDelayType                   := 0 ns;
--            tsetup_CLOCK_ENABLE_OUTPUT_CLK_posedge_posedge   : VitalDelayType                   := 0 ns;
--			tsetup_D_OUT_0_OUTPUT_CLK_negedge_posedge   : VitalDelayType                   := 0 ns;
--            tsetup_D_OUT_0_OUTPUT_CLK_posedge_posedge   : VitalDelayType                   := 0 ns;
--			tsetup_D_OUT_1_OUTPUT_CLK_negedge_negedge   : VitalDelayType                   := 0 ns;
--            tsetup_D_OUT_1_OUTPUT_CLK_posedge_negedge   : VitalDelayType                   := 0 ns;
--			tsetup_OUTPUT_ENABLE_OUTPUT_CLK_negedge_posedge   : VitalDelayType                   := 0 ns;
--            tsetup_OUTPUT_ENABLE_OUTPUT_CLK_posedge_posedge   : VitalDelayType                   := 0 ns;
--			--- VITAL hold time 
--			thold_CLOCK_ENABLE_INPUT_CLK_negedge_posedge    : VitalDelayType                   := 0 ns;
--            thold_CLOCK_ENABLE_INPUT_CLK_posedge_posedge    : VitalDelayType                   := 0 ns;
--            thold_PACKAGE_PIN_INPUT_CLK_negedge_posedge : VitalDelayType                   := 0 ns;
--            thold_PACKAGE_PIN_INPUT_CLK_posedge_posedge : VitalDelayType                   := 0 ns;
--            thold_PACKAGE_PIN_INPUT_CLK_posedge_negedge : VitalDelayType                   := 0 ns;
--            thold_PACKAGE_PIN_INPUT_CLK_negedge_negedge : VitalDelayType                   := 0 ns;
--            thold_CLOCK_ENABLE_OUTPUT_CLK_negedge_posedge   : VitalDelayType                   := 0 ns;
--            thold_CLOCK_ENABLE_OUTPUT_CLK_posedge_posedge   : VitalDelayType                   := 0 ns;
--			thold_D_OUT_0_OUTPUT_CLK_negedge_posedge   : VitalDelayType                   := 0 ns;
--            thold_D_OUT_0_OUTPUT_CLK_posedge_posedge   : VitalDelayType                   := 0 ns;
--			thold_D_OUT_1_OUTPUT_CLK_negedge_negedge   : VitalDelayType                   := 0 ns;
--            thold_D_OUT_1_OUTPUT_CLK_posedge_negedge   : VitalDelayType                   := 0 ns;
--			thold_OUTPUT_ENABLE_OUTPUT_CLK_negedge_posedge   : VitalDelayType                   := 0 ns;
--            thold_OUTPUT_ENABLE_OUTPUT_CLK_posedge_posedge   : VitalDelayType                   := 0 ns
--			
-- 			);
--	port 
--		(
--		D_OUT_1 		    : in std_logic;
--		D_OUT_0 		    : in std_logic;
--		CLOCK_ENABLE		: in std_logic;
--		LATCH_INPUT_VALUE	: in std_logic;
--		INPUT_CLK			: in std_logic;
--		
--		D_IN_1				: out std_logic;
--		D_IN_0				: out std_logic;
--		OUTPUT_ENABLE		: in std_logic;
--		OUTPUT_CLK			: in std_logic;
--		PACKAGE_PIN			: inout	std_logic
--		); 
--	attribute VITAL_LEVEL0 of
--      SB_IO : entity is true;	
--end SB_IO ;
--
--architecture SB_IO_V of SB_IO is
--  attribute VITAL_LEVEL0 of
--    SB_IO_V : architecture is true;
--
--	component	preio_physical
--	port	(
--			hold	:	in 	std_logic;
--			rstio	:	in	std_logic;
--			bs_en	:	in	std_logic;
--			shift	:	in	std_logic;
--			tclk	:	in	std_logic;
--			inclk	:	in	std_logic;
--			outclk	:	in	std_logic;
--			update	:	in	std_logic;
--			oepin	:	in	std_logic;
--			sdi		:	in	std_logic;
--			mode	:	in	std_logic;
--			hiz_b	:	in	std_logic;
--			sdo		:	out	std_logic;
--			dout1	:	out	std_logic;
--			dout0	:	out	std_logic;
--			ddr1	:	in	std_logic;
--			ddr0	:	in	std_logic;
--			padin	:	in	std_logic;
--			padout	:	out	std_logic;
--			padoen	:	out	std_logic;
--			cbit	:	in	std_logic_vector	(5 downto 0)
--			);
--	end component;
--
--	
--	signal D_OUT_1_ipd : std_ulogic := 'X';
--    signal D_OUT_0_ipd  : std_ulogic := 'X';
--    signal CLOCK_ENABLE_ipd  : std_ulogic := 'X';
--    signal LATCH_INPUT_VALUE_ipd   : std_ulogic := 'X';
--	signal INPUT_CLK_ipd : std_ulogic := 'X';
--    signal OUTPUT_ENABLE_ipd  : std_ulogic := 'X';
--    signal OUTPUT_CLK_ipd  : std_ulogic := 'X';
--	signal PACKAGE_PIN_ipd : std_ulogic;   --input direction
--	
--	signal Violation : std_ulogic;
--	--signal PACKAGE_PIN_zd : std_ulogic;
--	signal D_IN_0_zd : std_ulogic;
--	signal D_IN_1_zd : std_ulogic;
--------------------------------------------------------------------------------------------------------------------------------------------------	
--	signal	inclk_n, outclk_n, inclk, outclk,sdo	:	std_logic;
--	
--	signal	bs_en	:	std_logic	:='0';	--Boundary scan enable           
--	signal	shift	:	std_logic	:='0';	--Boundary scan shift            
--	signal	tclk	:	std_logic	:='0';	--Boundary scan clock            
--	signal	update	:	std_logic	:='0';	--Boundary scan update           
--	signal	sdi		:	std_logic	:='0';	--Boundary scan serial data in   
--	signal	mode	:	std_logic	:='0';	--Boundary scan mode             
--	signal	hiz_b	:	std_logic	:='1';	--Boundary scan Tristate control 
--	
--	signal	pin_cbit:	std_logic_vector(5 downto 0);
--	signal	neg_trig:	std_logic;
--	signal	pull_up	:	std_logic;
--	
--	signal	hold,oepin,padoen,padout,padin	:	std_logic;	
------------------------------------------------------------------------------------------------------------------------------------------------------	
--begin
--      WireDelay   : block
--        begin
--          VitalWireDelay (D_OUT_1_ipd, D_OUT_1, tipd_D_OUT_1);
--          VitalWireDelay (D_OUT_0_ipd, D_OUT_0, tipd_D_OUT_0);
--          VitalWireDelay (CLOCK_ENABLE_ipd, CLOCK_ENABLE, tipd_CLOCK_ENABLE);
--          VitalWireDelay (LATCH_INPUT_VALUE_ipd, LATCH_INPUT_VALUE, tipd_LATCH_INPUT_VALUE);
--		  VitalWireDelay (INPUT_CLK_ipd, INPUT_CLK, tipd_INPUT_CLK);
--          VitalWireDelay (OUTPUT_ENABLE_ipd, OUTPUT_ENABLE, tipd_OUTPUT_ENABLE);
--          VitalWireDelay (OUTPUT_CLK_ipd, OUTPUT_CLK, tipd_OUTPUT_CLK);
--		  VitalWireDelay (PACKAGE_PIN_ipd, PACKAGE_PIN, tipd_PACKAGE_PIN);
--        end block;
--		
--
---------------------------------------------------------------------------------
---- BEHAVIOR SECTION
---------------------------------------------------------------------------------
--	pin_cbit	<=	TO_STDLOGICVECTOR	(PIN_TYPE);
--	neg_trig	<=	TO_STDLOGIC	(NEG_TRIGGER);
--	pull_up		<=	TO_STDLOGIC	(PULLUP);
--	
----	OUTPUT_ENABLE	<=	'H';		--	weak 1 for initial value
--	inclk_n	<= 	INPUT_CLK_ipd xor neg_trig;
--	outclk_n	<=	OUTPUT_CLK_ipd xor neg_trig;
--	inclk	<=	inclk_n and CLOCK_ENABLE_ipd;
--	outclk	<=	outclk_n and CLOCK_ENABLE_ipd;
--	
--	hold	<=	LATCH_INPUT_VALUE_ipd;
--	oepin	<=	OUTPUT_ENABLE_ipd;
--	
--	padin	<=	PACKAGE_PIN_ipd;
--	-----------------------------------------------------------------	
--	preio_physical_i	:	preio_physical
--	port map	(
--				hold	=>	hold,
--				rstio	=>	'0',
--				bs_en	=>	bs_en,
--				shift	=>	shift,
--				tclk	=>	tclk,
--				inclk	=>	inclk,
--				outclk	=>	outclk,
--				update	=>	update,
--				oepin	=>	oepin,
--				sdi		=>	sdi,
--				mode	=>	mode,
--				hiz_b	=>	hiz_b,
--				sdo		=>	sdo,
--				dout1	=>	D_IN_1_zd,
--				dout0	=>	D_IN_0_zd,
--				ddr1	=>	D_OUT_1,
--				ddr0	=>	D_OUT_0,
--				padin	=>	padin,
--				padout	=>	padout,
--				padoen	=>	padoen,
--				cbit	=>	pin_cbit
--				);
---------------------------------------------------------------------
----VITAL timing check
--------------------------------------------------------------------
--  VITALTimingCheck : process (D_OUT_1_ipd, D_OUT_0_ipd, CLOCK_ENABLE_ipd, LATCH_INPUT_VALUE_ipd, INPUT_CLK_ipd, OUTPUT_ENABLE_ipd, OUTPUT_CLK_ipd, PACKAGE_PIN_ipd)
--    variable Tviol_D_OUT_0_OUTPUT_CLK_posedge : std_ulogic := '0';
--    variable Tviol_OUTPUT_ENABLE_OUTPUT_CLK_posedge : std_ulogic := '0';
--    variable Tviol_CLOCK_ENABLE_OUTPUT_CLK_posedge : std_ulogic := '0';
--    variable Tviol_D_OUT_1_OUTPUT_CLK_negedge : std_ulogic := '0';
--    variable Tviol_CLOCK_ENABLE_INPUT_CLK_posedge    : std_ulogic := '0';
--    variable Tviol_PACKAGE_PIN_INPUT_CLK_posedge   : std_ulogic := '0';
--	variable Tviol_PACKAGE_PIN_INPUT_CLK_negedge   : std_ulogic := '0';
--
--    variable Tmkr_D_OUT_0_OUTPUT_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
--    variable Tmkr_OUTPUT_ENABLE_OUTPUT_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
--    variable Tmkr_CLOCK_ENABLE_OUTPUT_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
--    variable Tmkr_D_OUT_1_OUTPUT_CLK_negedge : VitalTimingDataType := VitalTimingDataInit;
--    variable Tmkr_CLOCK_ENABLE_INPUT_CLK_posedge    : VitalTimingDataType := VitalTimingDataInit;
--    variable Tmkr_PACKAGE_PIN_INPUT_CLK_posedge   : VitalTimingDataType := VitalTimingDataInit;
--	variable Tmkr_PACKAGE_PIN_INPUT_CLK_negedge   : VitalTimingDataType := VitalTimingDataInit;
--	
--	
--  begin
--    
--    if (TimingChecksOn) then
--      VitalSetupHoldCheck (
--        Violation      => Tviol_D_OUT_0_OUTPUT_CLK_posedge,
--        TimingData     => Tmkr_D_OUT_0_OUTPUT_CLK_posedge,
--        TestSignal     => D_OUT_0_ipd,
--        TestSignalName => "D_OUT_0",
--        RefSignal      => OUTPUT_CLK_ipd,
--        RefSignalName  => "OUTPUT_CLK",
--        SetupHigh      => tsetup_D_OUT_0_OUTPUT_CLK_posedge_posedge,
--        SetupLow       => tsetup_D_OUT_0_OUTPUT_CLK_negedge_posedge,
--        HoldLow        => thold_D_OUT_0_OUTPUT_CLK_negedge_posedge,
--        HoldHigh       => thold_D_OUT_0_OUTPUT_CLK_posedge_posedge,
--        CheckEnabled   => true,
--        RefTransition  => 'R',
--        HeaderMsg      => "/SB_IO",
--        Xon            => Xon,
--        MsgOn          => true,
--        MsgSeverity    => warning);
--	  
--	  VitalSetupHoldCheck (
--        Violation      => Tviol_OUTPUT_ENABLE_OUTPUT_CLK_posedge,
--        TimingData     => Tmkr_OUTPUT_ENABLE_OUTPUT_CLK_posedge,
--        TestSignal     => OUTPUT_ENABLE_ipd,
--        TestSignalName => "OUTPUT_ENABLE",
--        RefSignal      => OUTPUT_CLK_ipd,
--        RefSignalName  => "OUTPUT_CLK",
--        SetupHigh      => tsetup_OUTPUT_ENABLE_OUTPUT_CLK_posedge_posedge,
--        SetupLow       => tsetup_OUTPUT_ENABLE_OUTPUT_CLK_negedge_posedge,
--        HoldLow        => thold_OUTPUT_ENABLE_OUTPUT_CLK_negedge_posedge,
--        HoldHigh       => thold_OUTPUT_ENABLE_OUTPUT_CLK_posedge_posedge,
--        CheckEnabled   => true,
--        RefTransition  => 'R',
--        HeaderMsg      => "/SB_IO",
--        Xon            => Xon,
--        MsgOn          => true,
--        MsgSeverity    => warning);
--		
--	  VitalSetupHoldCheck (
--        Violation      => Tviol_CLOCK_ENABLE_OUTPUT_CLK_posedge,
--        TimingData     => Tmkr_CLOCK_ENABLE_OUTPUT_CLK_posedge,
--        TestSignal     => CLOCK_ENABLE_ipd,
--        TestSignalName => "CLOCK_ENABLE",
--        RefSignal      => OUTPUT_CLK_ipd,
--        RefSignalName  => "OUTPUT_CLK",
--        SetupHigh      => tsetup_CLOCK_ENABLE_OUTPUT_CLK_posedge_posedge,
--        SetupLow       => tsetup_CLOCK_ENABLE_OUTPUT_CLK_negedge_posedge,
--        HoldLow        => thold_CLOCK_ENABLE_OUTPUT_CLK_negedge_posedge,
--        HoldHigh       => thold_CLOCK_ENABLE_OUTPUT_CLK_posedge_posedge,
--        CheckEnabled   => true,
--        RefTransition  => 'R',
--        HeaderMsg      => "/SB_IO",
--        Xon            => Xon,
--        MsgOn          => true,
--        MsgSeverity    => warning);
--		
--	  VitalSetupHoldCheck (
--        Violation      => Tviol_D_OUT_1_OUTPUT_CLK_negedge,
--        TimingData     => Tmkr_D_OUT_1_OUTPUT_CLK_negedge,
--        TestSignal     => D_OUT_1_ipd,
--        TestSignalName => "D_OUT_1",
--        RefSignal      => OUTPUT_CLK_ipd,
--        RefSignalName  => "OUTPUT_CLK",
--        SetupHigh      => tsetup_D_OUT_1_OUTPUT_CLK_negedge_negedge,
--        SetupLow       => tsetup_D_OUT_1_OUTPUT_CLK_posedge_negedge,
--        HoldLow        => thold_D_OUT_1_OUTPUT_CLK_negedge_negedge,
--        HoldHigh       => thold_D_OUT_1_OUTPUT_CLK_posedge_negedge,
--        CheckEnabled   => true,
--        RefTransition  => 'R',
--        HeaderMsg      => "/SB_IO",
--        Xon            => Xon,
--        MsgOn          => true,
--        MsgSeverity    => warning);
--		
--      VitalSetupHoldCheck (
--        Violation      => Tviol_CLOCK_ENABLE_INPUT_CLK_posedge,
--        TimingData     => Tmkr_CLOCK_ENABLE_INPUT_CLK_posedge,
--        TestSignal     => CLOCK_ENABLE_ipd,
--        TestSignalName => "CLOCK_ENABLE",
--        RefSignal      => INPUT_CLK_ipd,
--        RefSignalName  => "INPUT_CLK",
--        SetupHigh      => tsetup_CLOCK_ENABLE_INPUT_CLK_posedge_posedge,
--        SetupLow       => tsetup_CLOCK_ENABLE_INPUT_CLK_negedge_posedge,
--        HoldLow        => thold_CLOCK_ENABLE_INPUT_CLK_negedge_posedge,
--        HoldHigh       => thold_CLOCK_ENABLE_INPUT_CLK_posedge_posedge,
--        CheckEnabled   => true,
--        RefTransition  => 'R',
--        HeaderMsg      => "/SB_IO",
--        Xon            => Xon,
--        MsgOn          => true,
--        MsgSeverity    => warning);
--	  VitalSetupHoldCheck (
--        Violation      => Tviol_PACKAGE_PIN_INPUT_CLK_posedge,
--        TimingData     => Tmkr_PACKAGE_PIN_INPUT_CLK_posedge,
--        TestSignal     => PACKAGE_PIN_ipd,
--        TestSignalName => "PACKAGE_PIN",
--        RefSignal      => INPUT_CLK_ipd,
--        RefSignalName  => "INPUT_CLK",
--        SetupHigh      => tsetup_PACKAGE_PIN_INPUT_CLK_posedge_posedge,
--        SetupLow       => tsetup_PACKAGE_PIN_INPUT_CLK_negedge_posedge,
--        HoldLow        => thold_PACKAGE_PIN_INPUT_CLK_negedge_posedge,
--        HoldHigh       => thold_PACKAGE_PIN_INPUT_CLK_posedge_posedge,
--        CheckEnabled   => true,
--        RefTransition  => 'R',
--        HeaderMsg      => "/SB_IO",
--        Xon            => Xon,
--        MsgOn          => true,
--        MsgSeverity    => warning);
--		
--	  VitalSetupHoldCheck (
--        Violation      => Tviol_PACKAGE_PIN_INPUT_CLK_negedge,
--        TimingData     => Tmkr_PACKAGE_PIN_INPUT_CLK_negedge,
--        TestSignal     => PACKAGE_PIN_ipd,
--        TestSignalName => "PACKAGE_PIN",
--        RefSignal      => INPUT_CLK_ipd,
--        RefSignalName  => "INPUT_CLK",
--        SetupHigh      => tsetup_PACKAGE_PIN_INPUT_CLK_negedge_negedge,
--        SetupLow       => tsetup_PACKAGE_PIN_INPUT_CLK_posedge_negedge,
--        HoldLow        => thold_PACKAGE_PIN_INPUT_CLK_negedge_negedge,
--        HoldHigh       => thold_PACKAGE_PIN_INPUT_CLK_posedge_negedge,
--        CheckEnabled   => true,
--        RefTransition  => 'R',
--        HeaderMsg      => "/SB_IO",
--        Xon            => Xon,
--        MsgOn          => true,
--        MsgSeverity    => warning);
--     
--    end if;
--end process VITALTimingCheck;
----path delay
--  VITALPathDelay          : process (padout, padoen, D_OUT_1_ipd, D_OUT_0_ipd, PACKAGE_PIN_ipd, CLOCK_ENABLE_ipd, OUTPUT_ENABLE_ipd, LATCH_INPUT_VALUE_ipd, D_IN_0_zd, D_IN_1_zd, OUTPUT_CLK_ipd, INPUT_CLK_ipd)
--    variable PACKAGE_PIN_GlitchData : VitalGlitchDataType;
--	variable D_IN_0_GlitchData : VitalGlitchDataType;
--	variable D_IN_1_GlitchData : VitalGlitchDataType;
--	
--	variable tmp_padio : std_logic;  --package_pin output direction
--
--  begin
--   -- padin	<=	PACKAGE_PIN_ipd;
--		if	(padoen='1') then
--			tmp_padio	:=	'Z';
--		else
--			tmp_padio	:=	padout;
--		end if;
--  VitalPathDelay01 (
--      OutSignal                 => PACKAGE_PIN,
--      GlitchData                => PACKAGE_PIN_GlitchData,
--      OutSignalName             => "PACKAGE_PIN",
--      OutTemp                   => tmp_padio,
--      Paths                     => (0 => (D_OUT_0_ipd'last_event, tpd_D_OUT_0_PACKAGE_PIN, true),
--                                    1 => (D_OUT_1_ipd'last_event, tpd_D_OUT_1_PACKAGE_PIN, true),
--									2 => (OUTPUT_ENABLE_ipd'last_event, tpd_OUTPUT_ENABLE_PACKAGE_PIN, true),
--									3 => (OUTPUT_CLK_ipd'last_event, tpd_OUTPUT_CLK_PACKAGE_PIN, true)
--									),
--      Mode                      => VitalTransport,
--      Xon                       => Xon,
--      MsgOn                     => MsgOn,
--      MsgSeverity               => warning);
--	  
--	VitalPathDelay01 (
--      OutSignal                 => D_IN_0,
--      GlitchData                => D_IN_0_GlitchData,
--      OutSignalName             => "D_IN_0",
--      OutTemp                   => D_IN_0_zd,
--      Paths                     => (0 => (LATCH_INPUT_VALUE_ipd'last_event, tpd_LATCH_INPUT_VALUE_D_IN_0, true),
--									1 => (INPUT_CLK_ipd'last_event, tpd_INPUT_CLK_D_IN_0, true),
--									2 => (PACKAGE_PIN_ipd'last_event, tpd_PACKAGE_PIN_D_IN_0, true)
--									),
--      Mode                      => VitalTransport,
--      Xon                       => Xon,
--      MsgOn                     => MsgOn,
--      MsgSeverity               => warning);
--	  
--	VitalPathDelay01 (
--      OutSignal                 => D_IN_1,
--      GlitchData                => D_IN_1_GlitchData,
--      OutSignalName             => "D_IN_1",
--      OutTemp                   => D_IN_1_zd,
--      Paths                     => (0 => (LATCH_INPUT_VALUE_ipd'last_event, tpd_LATCH_INPUT_VALUE_D_IN_1, true),
--									1 => (INPUT_CLK_ipd'last_event, tpd_INPUT_CLK_D_IN_1, true),
--									2 => (PACKAGE_PIN_ipd'last_event, tpd_PACKAGE_PIN_D_IN_1, true)
--									),
--      Mode                      => VitalTransport,
--      Xon                       => Xon,
--      MsgOn                     => MsgOn,
--      MsgSeverity               => warning);
--  end process VITALPathDelay;
--
--
--end	SB_IO_V;

----------------------------------------------------------------------
--					SB_GB_IO
----------------------------------------------------------------------
--library ieee;
--use ieee.std_logic_1164.all;
--use ieee.std_logic_arith.all;
--use ieee.std_logic_unsigned.all;
--use IEEE.Vital_Primitives.all;
--use IEEE.VITAL_Timing.all;
----library	work;
--use	work.std_logic_SBT.all;
--
--entity	SB_GB_IO is
--	generic (
--			NEG_TRIGGER : bit						:=	'0';
--			PIN_TYPE	: bit_vector (5 downto 0)	:=	"000000";
--			PULLUP		: bit						:=	'0';
--			IO_STANDARD	: string					:=	"SB_LVCMOS";
--			----------------------------------------------------------------------------------
--			--VITAL PARAMETER
--			---------------------------------------------------------------------------------
--			TimingChecksOn  : boolean := true;
--			Xon   : boolean := true;
--            MsgOn : boolean := false;
--			--- VITAL path delay
--			tipd_D_OUT_1       : VitalDelayType01 := (0 ns, 0 ns);
--            tipd_D_OUT_0       : VitalDelayType01 := (0 ns, 0 ns);
--            tipd_CLOCK_ENABLE        : VitalDelayType01 := (0 ns, 0 ns);
--            tipd_LATCH_INPUT_VALUE       : VitalDelayType01 := (0 ns, 0 ns);
--            tipd_INPUT_CLK        : VitalDelayType01 := (0 ns, 0 ns);
--			tipd_OUTPUT_ENABLE       : VitalDelayType01 := (0 ns, 0 ns);
--            tipd_OUTPUT_CLK       : VitalDelayType01 := (0 ns, 0 ns);
--			tipd_PACKAGE_PIN      : VitalDelayType01 := (0 ns, 0 ns);
--            --- VITAL path delay
--            tpd_PACKAGE_PIN_D_IN_0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
--            tpd_PACKAGE_PIN_D_IN_1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
--            tpd_D_OUT_0_PACKAGE_PIN : VitalDelayType01 := (0.000 ns, 0.000 ns);
--			tpd_D_OUT_1_PACKAGE_PIN : VitalDelayType01 := (0.000 ns, 0.000 ns);
--            tpd_OUTPUT_ENABLE_PACKAGE_PIN : VitalDelayType01 := (0.000 ns, 0.000 ns);
--            tpd_LATCH_INPUT_VALUE_D_IN_0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
--			tpd_LATCH_INPUT_VALUE_D_IN_1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
--			tpd_PACKAGE_PIN_GLOBAL_BUFFER_OUTPUT : VitalDelayType01 := (0.000 ns, 0.000 ns);
--			--  VITAL clk-to-output path delay
--			tpd_INPUT_CLK_D_IN_0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
--            tpd_INPUT_CLK_D_IN_1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
--			tpd_OUTPUT_CLK_PACKAGE_PIN : VitalDelayType01 := (0.000 ns, 0.000 ns);
--			--- VITAL setup time
--			tsetup_CLOCK_ENABLE_INPUT_CLK_negedge_posedge    : VitalDelayType                   := 0 ns;
--            tsetup_CLOCK_ENABLE_INPUT_CLK_posedge_posedge    : VitalDelayType                   := 0 ns;
--            tsetup_PACKAGE_PIN_INPUT_CLK_negedge_posedge : VitalDelayType                   := 0 ns;
--            tsetup_PACKAGE_PIN_INPUT_CLK_posedge_posedge : VitalDelayType                   := 0 ns;
--            tsetup_PACKAGE_PIN_INPUT_CLK_posedge_negedge : VitalDelayType                   := 0 ns;
--            tsetup_PACKAGE_PIN_INPUT_CLK_negedge_negedge : VitalDelayType                   := 0 ns;
--            tsetup_CLOCK_ENABLE_OUTPUT_CLK_negedge_posedge   : VitalDelayType                   := 0 ns;
--            tsetup_CLOCK_ENABLE_OUTPUT_CLK_posedge_posedge   : VitalDelayType                   := 0 ns;
--			tsetup_D_OUT_0_OUTPUT_CLK_negedge_posedge   : VitalDelayType                   := 0 ns;
--            tsetup_D_OUT_0_OUTPUT_CLK_posedge_posedge   : VitalDelayType                   := 0 ns;
--			tsetup_D_OUT_1_OUTPUT_CLK_negedge_negedge   : VitalDelayType                   := 0 ns;
--            tsetup_D_OUT_1_OUTPUT_CLK_posedge_negedge   : VitalDelayType                   := 0 ns;
--			tsetup_OUTPUT_ENABLE_OUTPUT_CLK_negedge_posedge   : VitalDelayType                   := 0 ns;
--            tsetup_OUTPUT_ENABLE_OUTPUT_CLK_posedge_posedge   : VitalDelayType                   := 0 ns;
--			--- VITAL hold time 
--			thold_CLOCK_ENABLE_INPUT_CLK_negedge_posedge    : VitalDelayType                   := 0 ns;
--            thold_CLOCK_ENABLE_INPUT_CLK_posedge_posedge    : VitalDelayType                   := 0 ns;
--            thold_PACKAGE_PIN_INPUT_CLK_negedge_posedge : VitalDelayType                   := 0 ns;
--            thold_PACKAGE_PIN_INPUT_CLK_posedge_posedge : VitalDelayType                   := 0 ns;
--            thold_PACKAGE_PIN_INPUT_CLK_posedge_negedge : VitalDelayType                   := 0 ns;
--            thold_PACKAGE_PIN_INPUT_CLK_negedge_negedge : VitalDelayType                   := 0 ns;
--            thold_CLOCK_ENABLE_OUTPUT_CLK_negedge_posedge   : VitalDelayType                   := 0 ns;
--            thold_CLOCK_ENABLE_OUTPUT_CLK_posedge_posedge   : VitalDelayType                   := 0 ns;
--			thold_D_OUT_0_OUTPUT_CLK_negedge_posedge   : VitalDelayType                   := 0 ns;
--            thold_D_OUT_0_OUTPUT_CLK_posedge_posedge   : VitalDelayType                   := 0 ns;
--			thold_D_OUT_1_OUTPUT_CLK_negedge_negedge   : VitalDelayType                   := 0 ns;
--            thold_D_OUT_1_OUTPUT_CLK_posedge_negedge   : VitalDelayType                   := 0 ns;
--			thold_OUTPUT_ENABLE_OUTPUT_CLK_negedge_posedge   : VitalDelayType                   := 0 ns;
--            thold_OUTPUT_ENABLE_OUTPUT_CLK_posedge_posedge   : VitalDelayType                   := 0 ns
--			
-- 			);
--			
--	port	(
--			PACKAGE_PIN			:	inout	std_logic;
--			LATCH_INPUT_VALUE	:	in		std_logic;
--			CLOCK_ENABLE        :	in		std_logic;
--			INPUT_CLK           :	in		std_logic;
--			OUTPUT_CLK          :	in		std_logic;
--			OUTPUT_ENABLE		: in std_logic	:='H';
--			D_OUT_1             :	in		std_logic;
--			D_OUT_0             :	in		std_logic;
--			D_IN_1              :	out		std_logic;
--			D_IN_0              :	out		std_logic;
--			GLOBAL_BUFFER_OUTPUT:	out		std_logic
--			);
--	attribute VITAL_LEVEL0 of
--      SB_GB_IO : entity is true;	
--end SB_GB_IO;
--
--architecture SB_GB_IO_V of SB_GB_IO is
--  attribute VITAL_LEVEL0 of
--    SB_GB_IO_V : architecture is true;
--
--	component	preio_physical
--	port	(
--			hold	:	in 	std_logic;
--			rstio	:	in	std_logic;
--			bs_en	:	in	std_logic;
--			shift	:	in	std_logic;
--			tclk	:	in	std_logic;
--			inclk	:	in	std_logic;
--			outclk	:	in	std_logic;
--			update	:	in	std_logic;
--			oepin	:	in	std_logic;
--			sdi		:	in	std_logic;
--			mode	:	in	std_logic;
--			hiz_b	:	in	std_logic;
--			sdo		:	out	std_logic;
--			dout1	:	out	std_logic;
--			dout0	:	out	std_logic;
--			ddr1	:	in	std_logic;
--			ddr0	:	in	std_logic;
--			padin	:	in	std_logic;
--			padout	:	out	std_logic;
--			padoen	:	out	std_logic;
--			cbit	:	in	std_logic_vector	(5 downto 0)
--			);
--	end component;
--	
--	signal D_OUT_1_ipd : std_ulogic := 'X';
--    signal D_OUT_0_ipd  : std_ulogic := 'X';
--    signal CLOCK_ENABLE_ipd  : std_ulogic := 'X';
--    signal LATCH_INPUT_VALUE_ipd   : std_ulogic := 'X';
--	signal INPUT_CLK_ipd : std_ulogic := 'X';
--    signal OUTPUT_ENABLE_ipd  : std_ulogic := 'X';
--    signal OUTPUT_CLK_ipd  : std_ulogic := 'X';
--	signal PACKAGE_PIN_ipd : std_ulogic;   --input direction
--	
--	signal Violation : std_ulogic;
--	--signal PACKAGE_PIN_zd : std_ulogic;
--	signal D_IN_0_zd : std_ulogic;
--	signal D_IN_1_zd : std_ulogic;
--	signal GLOBAL_BUFFER_OUTPUT_zd : std_ulogic;
--------------------------------------------------------------------------------------------------------------------------------------------------	
--	signal	inclk_n, outclk_n, inclk, outclk,sdo	:	std_logic;
--	
--	signal	bs_en	:	std_logic	:='0';	--Boundary scan enable           
--	signal	shift	:	std_logic	:='0';	--Boundary scan shift            
--	signal	tclk	:	std_logic	:='0';	--Boundary scan clock            
--	signal	update	:	std_logic	:='0';	--Boundary scan update           
--	signal	sdi		:	std_logic	:='0';	--Boundary scan serial data in   
--	signal	mode	:	std_logic	:='0';	--Boundary scan mode             
--	signal	hiz_b	:	std_logic	:='1';	--Boundary scan Tristate control 
--	
--	signal	pin_cbit:	std_logic_vector(5 downto 0);
--	signal	neg_trig:	std_logic;
--	signal	pull_up	:	std_logic;
--	
--	signal	hold,oepin,padoen,padout,padin	:	std_logic;	
------------------------------------------------------------------------------------------------------------------------------------------------------	
--begin
--      WireDelay   : block
--        begin
--          VitalWireDelay (D_OUT_1_ipd, D_OUT_1, tipd_D_OUT_1);
--          VitalWireDelay (D_OUT_0_ipd, D_OUT_0, tipd_D_OUT_0);
--          VitalWireDelay (CLOCK_ENABLE_ipd, CLOCK_ENABLE, tipd_CLOCK_ENABLE);
--          VitalWireDelay (LATCH_INPUT_VALUE_ipd, LATCH_INPUT_VALUE, tipd_LATCH_INPUT_VALUE);
--		  VitalWireDelay (INPUT_CLK_ipd, INPUT_CLK, tipd_INPUT_CLK);
--          VitalWireDelay (OUTPUT_ENABLE_ipd, OUTPUT_ENABLE, tipd_OUTPUT_ENABLE);
--          VitalWireDelay (OUTPUT_CLK_ipd, OUTPUT_CLK, tipd_OUTPUT_CLK);
--		  VitalWireDelay (PACKAGE_PIN_ipd, PACKAGE_PIN, tipd_PACKAGE_PIN);
--        end block;
--		
--
--		
--
---------------------------------------------------------------------------------
---- BEHAVIOR SECTION
---------------------------------------------------------------------------------
--	pin_cbit	<=	TO_STDLOGICVECTOR	(PIN_TYPE);
--	neg_trig	<=	TO_STDLOGIC	(NEG_TRIGGER);
--	pull_up		<=	TO_STDLOGIC	(PULLUP);
----	OUTPUT_ENABLE	<=	'H';		--	weak 1 for initial value
--	inclk_n	<= 	INPUT_CLK_ipd xor neg_trig;
--	outclk_n	<=	OUTPUT_CLK_ipd xor neg_trig;
--	inclk	<=	inclk_n and CLOCK_ENABLE_ipd;
--	outclk	<=	outclk_n and CLOCK_ENABLE_ipd;
--	
--	hold	<=	LATCH_INPUT_VALUE_ipd;
--	oepin	<=	OUTPUT_ENABLE_ipd;
--	padin	<=	PACKAGE_PIN_ipd;
--	GLOBAL_BUFFER_OUTPUT_zd	<=	padin;
-------------------------------------------------------------------	
--
--	preio_physical_i	:	preio_physical
--	port map	(
--				hold	=>	hold,
--				rstio	=>	'0',
--				bs_en	=>	bs_en,
--				shift	=>	shift,
--				tclk	=>	tclk,
--				inclk	=>	inclk,
--				outclk	=>	outclk,
--				update	=>	update,
--				oepin	=>	oepin,
--				sdi		=>	sdi,
--				mode	=>	mode,
--				hiz_b	=>	hiz_b,
--				sdo		=>	sdo,
--				dout1	=>	D_IN_1,
--				dout0	=>	D_IN_0,
--				ddr1	=>	D_OUT_1,
--				ddr0	=>	D_OUT_0,
--				padin	=>	padin,
--				padout	=>	padout,
--				padoen	=>	padoen,
--				cbit	=>	pin_cbit
--				);
--
---------------------------------------------------------------------
----VITAL timing check
--------------------------------------------------------------------
--  VITALTimingCheck : process (D_OUT_1_ipd, D_OUT_0_ipd, CLOCK_ENABLE_ipd, LATCH_INPUT_VALUE_ipd, INPUT_CLK_ipd, OUTPUT_ENABLE_ipd, OUTPUT_CLK_ipd, PACKAGE_PIN_ipd)
--    variable Tviol_D_OUT_0_OUTPUT_CLK_posedge : std_ulogic := '0';
--    variable Tviol_OUTPUT_ENABLE_OUTPUT_CLK_posedge : std_ulogic := '0';
--    variable Tviol_CLOCK_ENABLE_OUTPUT_CLK_posedge : std_ulogic := '0';
--    variable Tviol_D_OUT_1_OUTPUT_CLK_negedge : std_ulogic := '0';
--    variable Tviol_CLOCK_ENABLE_INPUT_CLK_posedge    : std_ulogic := '0';
--    variable Tviol_PACKAGE_PIN_INPUT_CLK_posedge   : std_ulogic := '0';
--	variable Tviol_PACKAGE_PIN_INPUT_CLK_negedge   : std_ulogic := '0';
--
--    variable Tmkr_D_OUT_0_OUTPUT_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
--    variable Tmkr_OUTPUT_ENABLE_OUTPUT_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
--    variable Tmkr_CLOCK_ENABLE_OUTPUT_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
--    variable Tmkr_D_OUT_1_OUTPUT_CLK_negedge : VitalTimingDataType := VitalTimingDataInit;
--    variable Tmkr_CLOCK_ENABLE_INPUT_CLK_posedge    : VitalTimingDataType := VitalTimingDataInit;
--    variable Tmkr_PACKAGE_PIN_INPUT_CLK_posedge   : VitalTimingDataType := VitalTimingDataInit;
--	variable Tmkr_PACKAGE_PIN_INPUT_CLK_negedge   : VitalTimingDataType := VitalTimingDataInit;
--	
--	
--  begin
--    
--    if (TimingChecksOn) then
--      VitalSetupHoldCheck (
--        Violation      => Tviol_D_OUT_0_OUTPUT_CLK_posedge,
--        TimingData     => Tmkr_D_OUT_0_OUTPUT_CLK_posedge,
--        TestSignal     => D_OUT_0_ipd,
--        TestSignalName => "D_OUT_0",
--        RefSignal      => OUTPUT_CLK_ipd,
--        RefSignalName  => "OUTPUT_CLK",
--        SetupHigh      => tsetup_D_OUT_0_OUTPUT_CLK_posedge_posedge,
--        SetupLow       => tsetup_D_OUT_0_OUTPUT_CLK_negedge_posedge,
--        HoldLow        => thold_D_OUT_0_OUTPUT_CLK_negedge_posedge,
--        HoldHigh       => thold_D_OUT_0_OUTPUT_CLK_posedge_posedge,
--        CheckEnabled   => true,
--        RefTransition  => 'R',
--        HeaderMsg      => "/SB_IO",
--        Xon            => Xon,
--        MsgOn          => true,
--        MsgSeverity    => warning);
--	  
--	  VitalSetupHoldCheck (
--        Violation      => Tviol_OUTPUT_ENABLE_OUTPUT_CLK_posedge,
--        TimingData     => Tmkr_OUTPUT_ENABLE_OUTPUT_CLK_posedge,
--        TestSignal     => OUTPUT_ENABLE_ipd,
--        TestSignalName => "OUTPUT_ENABLE",
--        RefSignal      => OUTPUT_CLK_ipd,
--        RefSignalName  => "OUTPUT_CLK",
--        SetupHigh      => tsetup_OUTPUT_ENABLE_OUTPUT_CLK_posedge_posedge,
--        SetupLow       => tsetup_OUTPUT_ENABLE_OUTPUT_CLK_negedge_posedge,
--        HoldLow        => thold_OUTPUT_ENABLE_OUTPUT_CLK_negedge_posedge,
--        HoldHigh       => thold_OUTPUT_ENABLE_OUTPUT_CLK_posedge_posedge,
--        CheckEnabled   => true,
--        RefTransition  => 'R',
--        HeaderMsg      => "/SB_IO",
--        Xon            => Xon,
--        MsgOn          => true,
--        MsgSeverity    => warning);
--		
--	  VitalSetupHoldCheck (
--        Violation      => Tviol_CLOCK_ENABLE_OUTPUT_CLK_posedge,
--        TimingData     => Tmkr_CLOCK_ENABLE_OUTPUT_CLK_posedge,
--        TestSignal     => CLOCK_ENABLE_ipd,
--        TestSignalName => "CLOCK_ENABLE",
--        RefSignal      => OUTPUT_CLK_ipd,
--        RefSignalName  => "OUTPUT_CLK",
--        SetupHigh      => tsetup_CLOCK_ENABLE_OUTPUT_CLK_posedge_posedge,
--        SetupLow       => tsetup_CLOCK_ENABLE_OUTPUT_CLK_negedge_posedge,
--        HoldLow        => thold_CLOCK_ENABLE_OUTPUT_CLK_negedge_posedge,
--        HoldHigh       => thold_CLOCK_ENABLE_OUTPUT_CLK_posedge_posedge,
--        CheckEnabled   => true,
--        RefTransition  => 'R',
--        HeaderMsg      => "/SB_IO",
--        Xon            => Xon,
--        MsgOn          => true,
--        MsgSeverity    => warning);
--		
--	  VitalSetupHoldCheck (
--        Violation      => Tviol_D_OUT_1_OUTPUT_CLK_negedge,
--        TimingData     => Tmkr_D_OUT_1_OUTPUT_CLK_negedge,
--        TestSignal     => D_OUT_1_ipd,
--        TestSignalName => "D_OUT_1",
--        RefSignal      => OUTPUT_CLK_ipd,
--        RefSignalName  => "OUTPUT_CLK",
--        SetupHigh      => tsetup_D_OUT_1_OUTPUT_CLK_negedge_negedge,
--        SetupLow       => tsetup_D_OUT_1_OUTPUT_CLK_posedge_negedge,
--        HoldLow        => thold_D_OUT_1_OUTPUT_CLK_negedge_negedge,
--        HoldHigh       => thold_D_OUT_1_OUTPUT_CLK_posedge_negedge,
--        CheckEnabled   => true,
--        RefTransition  => 'R',
--        HeaderMsg      => "/SB_IO",
--        Xon            => Xon,
--        MsgOn          => true,
--        MsgSeverity    => warning);
--		
--      VitalSetupHoldCheck (
--        Violation      => Tviol_CLOCK_ENABLE_INPUT_CLK_posedge,
--        TimingData     => Tmkr_CLOCK_ENABLE_INPUT_CLK_posedge,
--        TestSignal     => CLOCK_ENABLE_ipd,
--        TestSignalName => "CLOCK_ENABLE",
--        RefSignal      => INPUT_CLK_ipd,
--        RefSignalName  => "INPUT_CLK",
--        SetupHigh      => tsetup_CLOCK_ENABLE_INPUT_CLK_posedge_posedge,
--        SetupLow       => tsetup_CLOCK_ENABLE_INPUT_CLK_negedge_posedge,
--        HoldLow        => thold_CLOCK_ENABLE_INPUT_CLK_negedge_posedge,
--        HoldHigh       => thold_CLOCK_ENABLE_INPUT_CLK_posedge_posedge,
--        CheckEnabled   => true,
--        RefTransition  => 'R',
--        HeaderMsg      => "/SB_IO",
--        Xon            => Xon,
--        MsgOn          => true,
--        MsgSeverity    => warning);
--	  VitalSetupHoldCheck (
--        Violation      => Tviol_PACKAGE_PIN_INPUT_CLK_posedge,
--        TimingData     => Tmkr_PACKAGE_PIN_INPUT_CLK_posedge,
--        TestSignal     => PACKAGE_PIN_ipd,
--        TestSignalName => "PACKAGE_PIN",
--        RefSignal      => INPUT_CLK_ipd,
--        RefSignalName  => "INPUT_CLK",
--        SetupHigh      => tsetup_PACKAGE_PIN_INPUT_CLK_posedge_posedge,
--        SetupLow       => tsetup_PACKAGE_PIN_INPUT_CLK_negedge_posedge,
--        HoldLow        => thold_PACKAGE_PIN_INPUT_CLK_negedge_posedge,
--        HoldHigh       => thold_PACKAGE_PIN_INPUT_CLK_posedge_posedge,
--        CheckEnabled   => true,
--        RefTransition  => 'R',
--        HeaderMsg      => "/SB_IO",
--        Xon            => Xon,
--        MsgOn          => true,
--        MsgSeverity    => warning);
--		
--	  VitalSetupHoldCheck (
--        Violation      => Tviol_PACKAGE_PIN_INPUT_CLK_negedge,
--        TimingData     => Tmkr_PACKAGE_PIN_INPUT_CLK_negedge,
--        TestSignal     => PACKAGE_PIN_ipd,
--        TestSignalName => "PACKAGE_PIN",
--        RefSignal      => INPUT_CLK_ipd,
--        RefSignalName  => "INPUT_CLK",
--        SetupHigh      => tsetup_PACKAGE_PIN_INPUT_CLK_negedge_negedge,
--        SetupLow       => tsetup_PACKAGE_PIN_INPUT_CLK_posedge_negedge,
--        HoldLow        => thold_PACKAGE_PIN_INPUT_CLK_negedge_negedge,
--        HoldHigh       => thold_PACKAGE_PIN_INPUT_CLK_posedge_negedge,
--        CheckEnabled   => true,
--        RefTransition  => 'R',
--        HeaderMsg      => "/SB_IO",
--        Xon            => Xon,
--        MsgOn          => true,
--        MsgSeverity    => warning);
--     
--    end if;
--end process VITALTimingCheck;
----path delay
--  VITALPathDelay          : process (padout, padoen, D_OUT_1_ipd, D_OUT_0_ipd, PACKAGE_PIN_ipd, CLOCK_ENABLE_ipd, OUTPUT_ENABLE_ipd, LATCH_INPUT_VALUE_ipd, D_IN_0_zd, D_IN_1_zd, GLOBAL_BUFFER_OUTPUT_zd)
--    variable PACKAGE_PIN_GlitchData : VitalGlitchDataType;
--	variable D_IN_0_GlitchData : VitalGlitchDataType;
--	variable D_IN_1_GlitchData : VitalGlitchDataType;
--	variable GLOBAL_BUFFER_OUTPUT_GlitchData : VitalGlitchDataType;
--	
--	variable tmp_padio : std_logic;  --package_pin output direction
--
--  begin
--    
--		if	(padoen='1') then
--			tmp_padio	:=	'Z';
--		else
--			tmp_padio	:=	padout;
--		end if;
--  VitalPathDelay01 (
--      OutSignal                 => PACKAGE_PIN,
--      GlitchData                => PACKAGE_PIN_GlitchData,
--      OutSignalName             => "PACKAGE_PIN",
--      OutTemp                   => tmp_padio,
--      Paths                     => (0 => (D_OUT_0_ipd'last_event, tpd_D_OUT_0_PACKAGE_PIN, true),
--                                    1 => (D_OUT_1_ipd'last_event, tpd_D_OUT_1_PACKAGE_PIN, true),
--									2 => (OUTPUT_ENABLE_ipd'last_event, tpd_OUTPUT_ENABLE_PACKAGE_PIN, true),
--									3 => (OUTPUT_CLK_ipd'last_event, tpd_OUTPUT_CLK_PACKAGE_PIN, true)
--									),
--      Mode                      => VitalTransport,
--      Xon                       => Xon,
--      MsgOn                     => MsgOn,
--      MsgSeverity               => warning);
--	  
--	VitalPathDelay01 (
--      OutSignal                 => D_IN_0,
--      GlitchData                => D_IN_0_GlitchData,
--      OutSignalName             => "D_IN_0",
--      OutTemp                   => D_IN_0_zd,
--      Paths                     => (0 => (LATCH_INPUT_VALUE_ipd'last_event, tpd_LATCH_INPUT_VALUE_D_IN_0, true),
--									1 => (INPUT_CLK_ipd'last_event, tpd_INPUT_CLK_D_IN_0, true),
--									2 => (PACKAGE_PIN_ipd'last_event, tpd_PACKAGE_PIN_D_IN_0, true)
--									),
--      Mode                      => VitalTransport,
--      Xon                       => Xon,
--      MsgOn                     => MsgOn,
--      MsgSeverity               => warning);
--	  
--	VitalPathDelay01 (
--      OutSignal                 => D_IN_1,
--      GlitchData                => D_IN_1_GlitchData,
--      OutSignalName             => "D_IN_1",
--      OutTemp                   => D_IN_1_zd,
--      Paths                     => (0 => (LATCH_INPUT_VALUE_ipd'last_event, tpd_LATCH_INPUT_VALUE_D_IN_1, true),
--									1 => (INPUT_CLK_ipd'last_event, tpd_INPUT_CLK_D_IN_1, true),
--									2 => (PACKAGE_PIN_ipd'last_event, tpd_PACKAGE_PIN_D_IN_1, true)
--									),
--      Mode                      => VitalTransport,
--      Xon                       => Xon,
--      MsgOn                     => MsgOn,
--      MsgSeverity               => warning);
--	  
--	VitalPathDelay01 (
--      OutSignal                 => GLOBAL_BUFFER_OUTPUT,
--      GlitchData                => GLOBAL_BUFFER_OUTPUT_GlitchData,
--      OutSignalName             => "GLOBAL_BUFFER_OUTPUT",
--      OutTemp                   => GLOBAL_BUFFER_OUTPUT_zd,
--      Paths                     => (0 => (PACKAGE_PIN_ipd'last_event, tpd_PACKAGE_PIN_D_IN_0, true)
--									),
--      Mode                      => VitalTransport,
--      Xon                       => Xon,
--      MsgOn                     => MsgOn,
--      MsgSeverity               => warning);
--  end process VITALPathDelay;
--end	SB_GB_IO_V;
--
-----------------------------------------------------------------
--					SB_GB
-----------------------------------------------------------------

--library ieee;
--use ieee.std_logic_1164.all;
--use ieee.std_logic_arith.all;
--use ieee.std_logic_unsigned.all;
--use IEEE.Vital_Primitives.all;
--use IEEE.VITAL_Timing.all;
----library	work;
--use	work.std_logic_SBT.all;
--
--entity	SB_GB	is
--generic	(----------------------------------------------------------------------------------
--			--VITAL PARAMETER
--			---------------------------------------------------------------------------------
--			TimingChecksOn  : boolean := true;
--			Xon   : boolean := true;
--            MsgOn : boolean := false;
--			--- VITAL path delay
--			tipd_USER_SIGNAL_TO_GLOBAL_BUFFER       : VitalDelayType01 := (0 ns, 0 ns);
--            --- VITAL path delay
--            tpd_USER_SIGNAL_TO_GLOBAL_BUFFER_GLOBAL_BUFFER_OUTPUT : VitalDelayType01 := (0.000 ns, 0.000 ns)
--            );
--port	(
--		GLOBAL_BUFFER_OUTPUT			:	out	std_logic;
--		USER_SIGNAL_TO_GLOBAL_BUFFER	:	in	std_logic
--		);
--attribute VITAL_LEVEL0 of
--      SB_GB : entity is true;
--end	SB_GB;
--
--architecture SB_GB_V of SB_GB is
--  attribute VITAL_LEVEL0 of
--    SB_GB_V : architecture is true;
--	
--  signal USER_SIGNAL_TO_GLOBAL_BUFFER_ipd   : std_ulogic := 'X';
--  signal GLOBAL_BUFFER_OUTPUT_zd : std_ulogic;
--  
--begin
--  WireDelay   : block
--        begin
--          VitalWireDelay (USER_SIGNAL_TO_GLOBAL_BUFFER_ipd, USER_SIGNAL_TO_GLOBAL_BUFFER, tipd_USER_SIGNAL_TO_GLOBAL_BUFFER);
--        end block;
----------------------------------------------------
----function part
---------------------------------------------------
--	GLOBAL_BUFFER_OUTPUT_zd	<=	USER_SIGNAL_TO_GLOBAL_BUFFER_ipd;
---------------------------------------------------------------------
----VITAL timing check
--------------------------------------------------------------------	
--	 VITALPathDelay          : process (USER_SIGNAL_TO_GLOBAL_BUFFER_ipd, GLOBAL_BUFFER_OUTPUT_zd)
-- --   variable O_zd         : std_ulogic;
--    variable O_GlitchData : VitalGlitchDataType;
--  begin
--    VitalPathDelay01 (
--      OutSignal                 => GLOBAL_BUFFER_OUTPUT,
--      GlitchData                => O_GlitchData,
--      OutSignalName             => "GLOBAL_BUFFER_OUTPUT",
--      OutTemp                   => GLOBAL_BUFFER_OUTPUT_zd,
--      Paths                     => (0 => (USER_SIGNAL_TO_GLOBAL_BUFFER_ipd'last_event, tpd_USER_SIGNAL_TO_GLOBAL_BUFFER_GLOBAL_BUFFER_OUTPUT, true)
-- 									),
--      Mode                      => VitalTransport,
--      Xon                       => Xon,
--      MsgOn                     => MsgOn,
--      MsgSeverity               => warning);
--  end process VITALPathDelay;
--end SB_GB_V;
--
--
--
--library ieee;
--use ieee.std_logic_1164.all;
--use ieee.std_logic_arith.all;
--use ieee.std_logic_unsigned.all;
--
--entity	SB_WARMBOOT	is
--port	(
--		BOOT	:	in	std_logic;
--		S1		:	in	std_logic;
--		S0		:	in	std_logic
--		);
--
--end SB_WARMBOOT;

-----------------------------------------------------------
--				SB_IO_DS
------------------------------------------------------------

--library ieee;
--use ieee.std_logic_1164.all;
--use ieee.std_logic_arith.all;
--use ieee.std_logic_unsigned.all;
--use IEEE.Vital_Primitives.all;
--use IEEE.VITAL_Timing.all;
----library	work;
--use	work.std_logic_SBT.all;
--
--entity	SB_IO_DS is
--	generic	(
--			NEG_TRIGGER : bit						:=	'0';
--			PIN_TYPE	: bit_vector (5 downto 0)	:=	"000000";
----			PULLUP		: bit						:=	'0';
--			IO_STANDARD	: string					:=	"SB_LVDS_OUTPUT";
--			----------------------------------------------------------------------------------
--			--VITAL PARAMETER
--			---------------------------------------------------------------------------------
--			TimingChecksOn  : boolean := true;
--			Xon   : boolean := true;
--            MsgOn : boolean := false;
--			--- VITAL path delay
--			tipd_D_OUT_1       : VitalDelayType01 := (0 ns, 0 ns);
--            tipd_D_OUT_0       : VitalDelayType01 := (0 ns, 0 ns);
--            tipd_CLOCK_ENABLE        : VitalDelayType01 := (0 ns, 0 ns);
--            tipd_LATCH_INPUT_VALUE       : VitalDelayType01 := (0 ns, 0 ns);
--            tipd_INPUT_CLK        : VitalDelayType01 := (0 ns, 0 ns);
--			tipd_OUTPUT_ENABLE       : VitalDelayType01 := (0 ns, 0 ns);
--            tipd_OUTPUT_CLK       : VitalDelayType01 := (0 ns, 0 ns);
--			tipd_PACKAGE_PIN      : VitalDelayType01 := (0 ns, 0 ns);
--            --- VITAL path delay
--            tpd_PACKAGE_PIN_D_IN_0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
--            tpd_PACKAGE_PIN_D_IN_1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
--            tpd_D_OUT_0_PACKAGE_PIN : VitalDelayType01 := (0.000 ns, 0.000 ns);
--			tpd_D_OUT_1_PACKAGE_PIN : VitalDelayType01 := (0.000 ns, 0.000 ns);
--            tpd_OUTPUT_ENABLE_PACKAGE_PIN : VitalDelayType01 := (0.000 ns, 0.000 ns);
--            tpd_LATCH_INPUT_VALUE_D_IN_0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
--			tpd_LATCH_INPUT_VALUE_D_IN_1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
--			tpd_D_OUT_0_PACKAGE_PIN_B : VitalDelayType01 := (0.000 ns, 0.000 ns);
--			tpd_D_OUT_1_PACKAGE_PIN_B : VitalDelayType01 := (0.000 ns, 0.000 ns);
--			tpd_OUTPUT_ENABLE_PACKAGE_PIN_B : VitalDelayType01 := (0.000 ns, 0.000 ns);
--			--  VITAL clk-to-output path delay
--			tpd_INPUT_CLK_D_IN_0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
--            tpd_INPUT_CLK_D_IN_1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
--			tpd_OUTPUT_CLK_PACKAGE_PIN : VitalDelayType01 := (0.000 ns, 0.000 ns);
--			tpd_OUTPUT_CLK_PACKAGE_PIN_B : VitalDelayType01 := (0.000 ns, 0.000 ns);
--			--- VITAL setup time
--			tsetup_CLOCK_ENABLE_INPUT_CLK_negedge_posedge    : VitalDelayType                   := 0 ns;
--            tsetup_CLOCK_ENABLE_INPUT_CLK_posedge_posedge    : VitalDelayType                   := 0 ns;
--            tsetup_PACKAGE_PIN_INPUT_CLK_negedge_posedge : VitalDelayType                   := 0 ns;
--            tsetup_PACKAGE_PIN_INPUT_CLK_posedge_posedge : VitalDelayType                   := 0 ns;
--            tsetup_PACKAGE_PIN_INPUT_CLK_posedge_negedge : VitalDelayType                   := 0 ns;
--            tsetup_PACKAGE_PIN_INPUT_CLK_negedge_negedge : VitalDelayType                   := 0 ns;
--            tsetup_CLOCK_ENABLE_OUTPUT_CLK_negedge_posedge   : VitalDelayType                   := 0 ns;
--            tsetup_CLOCK_ENABLE_OUTPUT_CLK_posedge_posedge   : VitalDelayType                   := 0 ns;
--			tsetup_D_OUT_0_OUTPUT_CLK_negedge_posedge   : VitalDelayType                   := 0 ns;
--            tsetup_D_OUT_0_OUTPUT_CLK_posedge_posedge   : VitalDelayType                   := 0 ns;
--			tsetup_D_OUT_1_OUTPUT_CLK_negedge_negedge   : VitalDelayType                   := 0 ns;
--            tsetup_D_OUT_1_OUTPUT_CLK_posedge_negedge   : VitalDelayType                   := 0 ns;
--			tsetup_OUTPUT_ENABLE_OUTPUT_CLK_negedge_posedge   : VitalDelayType                   := 0 ns;
--            tsetup_OUTPUT_ENABLE_OUTPUT_CLK_posedge_posedge   : VitalDelayType                   := 0 ns;
--			--- VITAL hold time 
--			thold_CLOCK_ENABLE_INPUT_CLK_negedge_posedge    : VitalDelayType                   := 0 ns;
--            thold_CLOCK_ENABLE_INPUT_CLK_posedge_posedge    : VitalDelayType                   := 0 ns;
--            thold_PACKAGE_PIN_INPUT_CLK_negedge_posedge : VitalDelayType                   := 0 ns;
--            thold_PACKAGE_PIN_INPUT_CLK_posedge_posedge : VitalDelayType                   := 0 ns;
--            thold_PACKAGE_PIN_INPUT_CLK_posedge_negedge : VitalDelayType                   := 0 ns;
--            thold_PACKAGE_PIN_INPUT_CLK_negedge_negedge : VitalDelayType                   := 0 ns;
--            thold_CLOCK_ENABLE_OUTPUT_CLK_negedge_posedge   : VitalDelayType                   := 0 ns;
--            thold_CLOCK_ENABLE_OUTPUT_CLK_posedge_posedge   : VitalDelayType                   := 0 ns;
--			thold_D_OUT_0_OUTPUT_CLK_negedge_posedge   : VitalDelayType                   := 0 ns;
--            thold_D_OUT_0_OUTPUT_CLK_posedge_posedge   : VitalDelayType                   := 0 ns;
--			thold_D_OUT_1_OUTPUT_CLK_negedge_negedge   : VitalDelayType                   := 0 ns;
--            thold_D_OUT_1_OUTPUT_CLK_posedge_negedge   : VitalDelayType                   := 0 ns;
--			thold_OUTPUT_ENABLE_OUTPUT_CLK_negedge_posedge   : VitalDelayType                   := 0 ns;
--            thold_OUTPUT_ENABLE_OUTPUT_CLK_posedge_posedge   : VitalDelayType                   := 0 ns
--			
--			);
--			
--	port	(
--			PACKAGE_PIN			:	inout	std_logic;
--			LATCH_INPUT_VALUE	:	in		std_logic;
--			CLOCK_ENABLE        :	in		std_logic;
--			INPUT_CLK           :	in		std_logic;
--			OUTPUT_CLK          :	in		std_logic;
--			OUTPUT_ENABLE		: in std_logic	:='H';
--			D_OUT_1             :	in		std_logic;
--			D_OUT_0             :	in		std_logic;
--			D_IN_1              :	out		std_logic;
--			D_IN_0              :	out		std_logic;
--			PACKAGE_PIN_B	    :	inout	std_logic	-- User's package pin - 'PAD' output  
--			);
--	attribute VITAL_LEVEL0 of
--      SB_IO_DS : entity is true;	
--end SB_IO_DS;
--
--architecture SB_IO_DS_V of SB_IO_DS is
--  attribute VITAL_LEVEL0 of
--    SB_IO_DS_V : architecture is true;
--
--	component	preio_physical
--	port	(
--			hold	:	in 	std_logic;
--			rstio	:	in	std_logic;
--			bs_en	:	in	std_logic;
--			shift	:	in	std_logic;
--			tclk	:	in	std_logic;
--			inclk	:	in	std_logic;
--			outclk	:	in	std_logic;
--			update	:	in	std_logic;
--			oepin	:	in	std_logic;
--			sdi		:	in	std_logic;
--			mode	:	in	std_logic;
--			hiz_b	:	in	std_logic;
--			sdo		:	out	std_logic;
--			dout1	:	out	std_logic;
--			dout0	:	out	std_logic;
--			ddr1	:	in	std_logic;
--			ddr0	:	in	std_logic;
--			padin	:	in	std_logic;
--			padout	:	out	std_logic;
--			padoen	:	out	std_logic;
--			cbit	:	in	std_logic_vector	(5 downto 0)
--			);
--	end component;
--	
--	signal D_OUT_1_ipd : std_ulogic := 'X';
--    signal D_OUT_0_ipd  : std_ulogic := 'X';
--    signal CLOCK_ENABLE_ipd  : std_ulogic := 'X';
--    signal LATCH_INPUT_VALUE_ipd   : std_ulogic := 'X';
--	signal INPUT_CLK_ipd : std_ulogic := 'X';
--    signal OUTPUT_ENABLE_ipd  : std_ulogic := 'X';
--    signal OUTPUT_CLK_ipd  : std_ulogic := 'X';
--	signal PACKAGE_PIN_ipd : std_ulogic;   --input direction
--	
--	signal Violation : std_ulogic;
--	--signal PACKAGE_PIN_zd : std_ulogic;
--	signal D_IN_0_zd : std_ulogic;
--	signal D_IN_1_zd : std_ulogic;
--------------------------------------------------------------------------------------------------------------------------------------------------	
--	signal	inclk_n, outclk_n, inclk, outclk,sdo	:	std_logic;
--	
--	signal	bs_en	:	std_logic	:='0';	--Boundary scan enable           
--	signal	shift	:	std_logic	:='0';	--Boundary scan shift            
--	signal	tclk	:	std_logic	:='0';	--Boundary scan clock            
--	signal	update	:	std_logic	:='0';	--Boundary scan update           
--	signal	sdi		:	std_logic	:='0';	--Boundary scan serial data in   
--	signal	mode	:	std_logic	:='0';	--Boundary scan mode             
--	signal	hiz_b	:	std_logic	:='1';	--Boundary scan Tristate control 
--	
--	signal	pin_cbit:	std_logic_vector(5 downto 0);
--	signal	neg_trig:	std_logic;
--	signal	pull_up	:	std_logic;
--	
--	signal	hold,oepin,padoen,padout,padin	:	std_logic;	
------------------------------------------------------------------------------------------------------------------------------------------------------	
--begin
--      WireDelay   : block
--        begin
--          VitalWireDelay (D_OUT_1_ipd, D_OUT_1, tipd_D_OUT_1);
--          VitalWireDelay (D_OUT_0_ipd, D_OUT_0, tipd_D_OUT_0);
--          VitalWireDelay (CLOCK_ENABLE_ipd, CLOCK_ENABLE, tipd_CLOCK_ENABLE);
--          VitalWireDelay (LATCH_INPUT_VALUE_ipd, LATCH_INPUT_VALUE, tipd_LATCH_INPUT_VALUE);
--		  VitalWireDelay (INPUT_CLK_ipd, INPUT_CLK, tipd_INPUT_CLK);
--          VitalWireDelay (OUTPUT_ENABLE_ipd, OUTPUT_ENABLE, tipd_OUTPUT_ENABLE);
--          VitalWireDelay (OUTPUT_CLK_ipd, OUTPUT_CLK, tipd_OUTPUT_CLK);
--		  VitalWireDelay (PACKAGE_PIN_ipd, PACKAGE_PIN, tipd_PACKAGE_PIN);
--        end block;
--		
--
---------------------------------------------------------------------------------
---- BEHAVIOR SECTION
---------------------------------------------------------------------------------
--	
--	pin_cbit	<=	TO_STDLOGICVECTOR	(PIN_TYPE);
--	neg_trig	<=	TO_STDLOGIC	(NEG_TRIGGER);
----	pull_up		<=	TO_STDLOGIC	(PULLUP);
--	
----	OUTPUT_ENABLE	<=	'H';		--	weak 1 for initial value
--	inclk_n	<= 	INPUT_CLK_ipd xor neg_trig;
--	outclk_n	<=	OUTPUT_CLK_ipd xor neg_trig;
--	inclk	<=	inclk_n and CLOCK_ENABLE_ipd;
--	outclk	<=	outclk_n and CLOCK_ENABLE_ipd;
--	
--	hold	<=	LATCH_INPUT_VALUE_ipd;
--	oepin	<=	OUTPUT_ENABLE_ipd;
--	
--	padin	<=	PACKAGE_PIN_ipd;
-------------------------------------------------------------------	
--
--	preio_physical_i	:	preio_physical
--	port map	(
--				hold	=>	hold,
--				rstio	=>	'0',
--				bs_en	=>	bs_en,
--				shift	=>	shift,
--				tclk	=>	tclk,
--				inclk	=>	inclk,
--				outclk	=>	outclk,
--				update	=>	update,
--				oepin	=>	oepin,
--				sdi		=>	sdi,
--				mode	=>	mode,
--				hiz_b	=>	hiz_b,
--				sdo		=>	sdo,
--				dout1	=>	D_IN_1,
--				dout0	=>	D_IN_0,
--				ddr1	=>	D_OUT_1,
--				ddr0	=>	D_OUT_0,
--				padin	=>	padin,
--				padout	=>	padout,
--				padoen	=>	padoen,
--				cbit	=>	pin_cbit
--				);
---------------------------------------------------------------------
----VITAL timing check
--------------------------------------------------------------------
--  VITALTimingCheck : process (D_OUT_1_ipd, D_OUT_0_ipd, CLOCK_ENABLE_ipd, LATCH_INPUT_VALUE_ipd, INPUT_CLK_ipd, OUTPUT_ENABLE_ipd, OUTPUT_CLK_ipd, PACKAGE_PIN_ipd)
--    variable Tviol_D_OUT_0_OUTPUT_CLK_posedge : std_ulogic := '0';
--    variable Tviol_OUTPUT_ENABLE_OUTPUT_CLK_posedge : std_ulogic := '0';
--    variable Tviol_CLOCK_ENABLE_OUTPUT_CLK_posedge : std_ulogic := '0';
--    variable Tviol_D_OUT_1_OUTPUT_CLK_negedge : std_ulogic := '0';
--    variable Tviol_CLOCK_ENABLE_INPUT_CLK_posedge    : std_ulogic := '0';
--    variable Tviol_PACKAGE_PIN_INPUT_CLK_posedge   : std_ulogic := '0';
--	variable Tviol_PACKAGE_PIN_INPUT_CLK_negedge   : std_ulogic := '0';
--
--    variable Tmkr_D_OUT_0_OUTPUT_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
--    variable Tmkr_OUTPUT_ENABLE_OUTPUT_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
--    variable Tmkr_CLOCK_ENABLE_OUTPUT_CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
--    variable Tmkr_D_OUT_1_OUTPUT_CLK_negedge : VitalTimingDataType := VitalTimingDataInit;
--    variable Tmkr_CLOCK_ENABLE_INPUT_CLK_posedge    : VitalTimingDataType := VitalTimingDataInit;
--    variable Tmkr_PACKAGE_PIN_INPUT_CLK_posedge   : VitalTimingDataType := VitalTimingDataInit;
--	variable Tmkr_PACKAGE_PIN_INPUT_CLK_negedge   : VitalTimingDataType := VitalTimingDataInit;
--	
--	
--  begin
--    
--    if (TimingChecksOn) then
--      VitalSetupHoldCheck (
--        Violation      => Tviol_D_OUT_0_OUTPUT_CLK_posedge,
--        TimingData     => Tmkr_D_OUT_0_OUTPUT_CLK_posedge,
--        TestSignal     => D_OUT_0_ipd,
--        TestSignalName => "D_OUT_0",
--        RefSignal      => OUTPUT_CLK_ipd,
--        RefSignalName  => "OUTPUT_CLK",
--        SetupHigh      => tsetup_D_OUT_0_OUTPUT_CLK_posedge_posedge,
--        SetupLow       => tsetup_D_OUT_0_OUTPUT_CLK_negedge_posedge,
--        HoldLow        => thold_D_OUT_0_OUTPUT_CLK_negedge_posedge,
--        HoldHigh       => thold_D_OUT_0_OUTPUT_CLK_posedge_posedge,
--        CheckEnabled   => true,
--        RefTransition  => 'R',
--        HeaderMsg      => "/SB_IO",
--        Xon            => Xon,
--        MsgOn          => true,
--        MsgSeverity    => warning);
--	  
--	  VitalSetupHoldCheck (
--        Violation      => Tviol_OUTPUT_ENABLE_OUTPUT_CLK_posedge,
--        TimingData     => Tmkr_OUTPUT_ENABLE_OUTPUT_CLK_posedge,
--        TestSignal     => OUTPUT_ENABLE_ipd,
--        TestSignalName => "OUTPUT_ENABLE",
--        RefSignal      => OUTPUT_CLK_ipd,
--        RefSignalName  => "OUTPUT_CLK",
--        SetupHigh      => tsetup_OUTPUT_ENABLE_OUTPUT_CLK_posedge_posedge,
--        SetupLow       => tsetup_OUTPUT_ENABLE_OUTPUT_CLK_negedge_posedge,
--        HoldLow        => thold_OUTPUT_ENABLE_OUTPUT_CLK_negedge_posedge,
--        HoldHigh       => thold_OUTPUT_ENABLE_OUTPUT_CLK_posedge_posedge,
--        CheckEnabled   => true,
--        RefTransition  => 'R',
--        HeaderMsg      => "/SB_IO",
--        Xon            => Xon,
--        MsgOn          => true,
--        MsgSeverity    => warning);
--		
--	  VitalSetupHoldCheck (
--        Violation      => Tviol_CLOCK_ENABLE_OUTPUT_CLK_posedge,
--        TimingData     => Tmkr_CLOCK_ENABLE_OUTPUT_CLK_posedge,
--        TestSignal     => CLOCK_ENABLE_ipd,
--        TestSignalName => "CLOCK_ENABLE",
--        RefSignal      => OUTPUT_CLK_ipd,
--        RefSignalName  => "OUTPUT_CLK",
--        SetupHigh      => tsetup_CLOCK_ENABLE_OUTPUT_CLK_posedge_posedge,
--        SetupLow       => tsetup_CLOCK_ENABLE_OUTPUT_CLK_negedge_posedge,
--        HoldLow        => thold_CLOCK_ENABLE_OUTPUT_CLK_negedge_posedge,
--        HoldHigh       => thold_CLOCK_ENABLE_OUTPUT_CLK_posedge_posedge,
--        CheckEnabled   => true,
--        RefTransition  => 'R',
--        HeaderMsg      => "/SB_IO",
--        Xon            => Xon,
--        MsgOn          => true,
--        MsgSeverity    => warning);
--		
--	  VitalSetupHoldCheck (
--        Violation      => Tviol_D_OUT_1_OUTPUT_CLK_negedge,
--        TimingData     => Tmkr_D_OUT_1_OUTPUT_CLK_negedge,
--        TestSignal     => D_OUT_1_ipd,
--        TestSignalName => "D_OUT_1",
--        RefSignal      => OUTPUT_CLK_ipd,
--        RefSignalName  => "OUTPUT_CLK",
--        SetupHigh      => tsetup_D_OUT_1_OUTPUT_CLK_negedge_negedge,
--        SetupLow       => tsetup_D_OUT_1_OUTPUT_CLK_posedge_negedge,
--        HoldLow        => thold_D_OUT_1_OUTPUT_CLK_negedge_negedge,
--        HoldHigh       => thold_D_OUT_1_OUTPUT_CLK_posedge_negedge,
--        CheckEnabled   => true,
--        RefTransition  => 'R',
--        HeaderMsg      => "/SB_IO",
--        Xon            => Xon,
--        MsgOn          => true,
--        MsgSeverity    => warning);
--		
--      VitalSetupHoldCheck (
--        Violation      => Tviol_CLOCK_ENABLE_INPUT_CLK_posedge,
--        TimingData     => Tmkr_CLOCK_ENABLE_INPUT_CLK_posedge,
--        TestSignal     => CLOCK_ENABLE_ipd,
--        TestSignalName => "CLOCK_ENABLE",
--        RefSignal      => INPUT_CLK_ipd,
--        RefSignalName  => "INPUT_CLK",
--        SetupHigh      => tsetup_CLOCK_ENABLE_INPUT_CLK_posedge_posedge,
--        SetupLow       => tsetup_CLOCK_ENABLE_INPUT_CLK_negedge_posedge,
--        HoldLow        => thold_CLOCK_ENABLE_INPUT_CLK_negedge_posedge,
--        HoldHigh       => thold_CLOCK_ENABLE_INPUT_CLK_posedge_posedge,
--        CheckEnabled   => true,
--        RefTransition  => 'R',
--        HeaderMsg      => "/SB_IO",
--        Xon            => Xon,
--        MsgOn          => true,
--        MsgSeverity    => warning);
--	  VitalSetupHoldCheck (
--        Violation      => Tviol_PACKAGE_PIN_INPUT_CLK_posedge,
--        TimingData     => Tmkr_PACKAGE_PIN_INPUT_CLK_posedge,
--        TestSignal     => PACKAGE_PIN_ipd,
--        TestSignalName => "PACKAGE_PIN",
--        RefSignal      => INPUT_CLK_ipd,
--        RefSignalName  => "INPUT_CLK",
--        SetupHigh      => tsetup_PACKAGE_PIN_INPUT_CLK_posedge_posedge,
--        SetupLow       => tsetup_PACKAGE_PIN_INPUT_CLK_negedge_posedge,
--        HoldLow        => thold_PACKAGE_PIN_INPUT_CLK_negedge_posedge,
--        HoldHigh       => thold_PACKAGE_PIN_INPUT_CLK_posedge_posedge,
--        CheckEnabled   => true,
--        RefTransition  => 'R',
--        HeaderMsg      => "/SB_IO",
--        Xon            => Xon,
--        MsgOn          => true,
--        MsgSeverity    => warning);
--		
--	  VitalSetupHoldCheck (
--        Violation      => Tviol_PACKAGE_PIN_INPUT_CLK_negedge,
--        TimingData     => Tmkr_PACKAGE_PIN_INPUT_CLK_negedge,
--        TestSignal     => PACKAGE_PIN_ipd,
--        TestSignalName => "PACKAGE_PIN",
--        RefSignal      => INPUT_CLK_ipd,
--        RefSignalName  => "INPUT_CLK",
--        SetupHigh      => tsetup_PACKAGE_PIN_INPUT_CLK_negedge_negedge,
--        SetupLow       => tsetup_PACKAGE_PIN_INPUT_CLK_posedge_negedge,
--        HoldLow        => thold_PACKAGE_PIN_INPUT_CLK_negedge_negedge,
--        HoldHigh       => thold_PACKAGE_PIN_INPUT_CLK_posedge_negedge,
--        CheckEnabled   => true,
--        RefTransition  => 'R',
--        HeaderMsg      => "/SB_IO",
--        Xon            => Xon,
--        MsgOn          => true,
--        MsgSeverity    => warning);
--     
--    end if;
--end process VITALTimingCheck;
----path delay
--  VITALPathDelay          : process (padout, padoen, D_OUT_1_ipd, D_OUT_0_ipd, PACKAGE_PIN_ipd, CLOCK_ENABLE_ipd, OUTPUT_ENABLE_ipd, LATCH_INPUT_VALUE_ipd, D_IN_0_zd, D_IN_1_zd, OUTPUT_CLK_ipd, INPUT_CLK_ipd)
--    variable PACKAGE_PIN_GlitchData : VitalGlitchDataType;
--	variable PACKAGE_PIN_B_GlitchData : VitalGlitchDataType;
--	variable D_IN_0_GlitchData : VitalGlitchDataType;
--	variable D_IN_1_GlitchData : VitalGlitchDataType;
--	
--	variable tmp_padio : std_logic;  --package_pin output direction
--	variable tmp_padio_b : std_logic;  --package_pin output direction
--
--  begin
-- 		if	(padoen='1') then
--			tmp_padio	:=	'Z';
--			tmp_padio_b	:=	'Z';
--		else
--			tmp_padio	:=	padout;
--			tmp_padio_b	:=	not padout;
--		end if;
--  VitalPathDelay01 (
--      OutSignal                 => PACKAGE_PIN,
--      GlitchData                => PACKAGE_PIN_GlitchData,
--      OutSignalName             => "PACKAGE_PIN",
--      OutTemp                   => tmp_padio,
--      Paths                     => (0 => (D_OUT_0_ipd'last_event, tpd_D_OUT_0_PACKAGE_PIN, true),
--                                    1 => (D_OUT_1_ipd'last_event, tpd_D_OUT_1_PACKAGE_PIN, true),
--									2 => (OUTPUT_ENABLE_ipd'last_event, tpd_OUTPUT_ENABLE_PACKAGE_PIN, true),
--									3 => (OUTPUT_CLK_ipd'last_event, tpd_OUTPUT_CLK_PACKAGE_PIN, true)
--									),
--      Mode                      => VitalTransport,
--      Xon                       => Xon,
--      MsgOn                     => MsgOn,
--      MsgSeverity               => warning);
--  VitalPathDelay01 (
--      OutSignal                 => PACKAGE_PIN_B,
--      GlitchData                => PACKAGE_PIN_B_GlitchData,
--      OutSignalName             => "PACKAGE_PIN_B",
--      OutTemp                   => tmp_padio_b,
--      Paths                     => (0 => (D_OUT_0_ipd'last_event, tpd_D_OUT_0_PACKAGE_PIN_B, true),
--                                    1 => (D_OUT_1_ipd'last_event, tpd_D_OUT_1_PACKAGE_PIN_B, true),
--									2 => (OUTPUT_ENABLE_ipd'last_event, tpd_OUTPUT_ENABLE_PACKAGE_PIN_B, true),
--									3 => (OUTPUT_CLK_ipd'last_event, tpd_OUTPUT_CLK_PACKAGE_PIN_B, true)
--									),
--      Mode                      => VitalTransport,
--      Xon                       => Xon,
--      MsgOn                     => MsgOn,
--      MsgSeverity               => warning);
--	  
--	VitalPathDelay01 (
--      OutSignal                 => D_IN_0,
--      GlitchData                => D_IN_0_GlitchData,
--      OutSignalName             => "D_IN_0",
--      OutTemp                   => D_IN_0_zd,
--      Paths                     => (0 => (LATCH_INPUT_VALUE_ipd'last_event, tpd_LATCH_INPUT_VALUE_D_IN_0, true),
--									1 => (INPUT_CLK_ipd'last_event, tpd_INPUT_CLK_D_IN_0, true),
--									2 => (PACKAGE_PIN_ipd'last_event, tpd_PACKAGE_PIN_D_IN_0, true)
--									),
--      Mode                      => VitalTransport,
--      Xon                       => Xon,
--      MsgOn                     => MsgOn,
--      MsgSeverity               => warning);
--	  
--	VitalPathDelay01 (
--      OutSignal                 => D_IN_1,
--      GlitchData                => D_IN_1_GlitchData,
--      OutSignalName             => "D_IN_1",
--      OutTemp                   => D_IN_1_zd,
--      Paths                     => (0 => (LATCH_INPUT_VALUE_ipd'last_event, tpd_LATCH_INPUT_VALUE_D_IN_1, true),
--									1 => (INPUT_CLK_ipd'last_event, tpd_INPUT_CLK_D_IN_1, true),
--									2 => (PACKAGE_PIN_ipd'last_event, tpd_PACKAGE_PIN_D_IN_1, true)
--									),
--      Mode                      => VitalTransport,
--      Xon                       => Xon,
--      MsgOn                     => MsgOn,
--      MsgSeverity               => warning);
--  end process VITALPathDelay;
--  
--end	SB_IO_DS_V;


-------------------------------------------------------------
--					GND
-------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity	GND	is
port	(
		Y	:	out	std_logic
		);

end GND;

architecture GND_V of GND is
begin
	Y	<=	'0';
end GND_V;

-------------------------------------------------------------
--					VCC
-------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity	VCC	is
port	(
		Y	:	out	std_logic
		);

end VCC;

architecture VCC_V of VCC is
begin
	Y	<=	'1';
end VCC_V;


----  Ligthning IP Primitives  ------- 

-----------------------------------------------
-----		  SB_I2C              	------- 
-----------------------------------------------
	
library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use IEEE.Vital_Primitives.all;
use IEEE.VITAL_Timing.all;
library WORK;
use WORK.vcomponent_vital.all;

entity  SB_I2C  is 
--define kinds of delay timing paras default value
	generic(
	I2C_SLAVE_INIT_ADDR : string := "0b1111100001";
	BUS_ADDR74 : string := "0b0001";
	-----------------------------------------------------------------
--VITAL PARAMETER	
	--------------------------------------------
TimingChecksOn  : boolean := true;
	Xon   : boolean := true;					   
    	MsgOn : boolean := false;
	--Vital path delay
Tipd_SBCLKI : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBRWI : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBSTBI : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBADRI7 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBADRI6 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBADRI5 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBADRI4 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBADRI3 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBADRI2 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBADRI1 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBADRI0 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBDATI7 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBDATI6 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBDATI5 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBDATI4 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBDATI3 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBDATI2 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBDATI1 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBDATI0 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SCLI : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SDAI : VitalDelayType01 := (0 ns, 0 ns);
--Tipd_SCLO : VitalDelayType01 := (0 ns, 0 ns);

--Vital path delay
tpd_SCLO_SDAO_posedge: VitalDelayType01 := (0.000 ns, 0.000 ns);	
tpd_SCLO_SDAOE_posedge: VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SCLI_SDAO_posedge: VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SCLI_SDAOE_posedge: VitalDelayType01 := (0.000 ns, 0.000 ns);
--Vital clk-to-output path delay
--tpd_SBCLKI_SCLO : VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SBCLKI_SBDATO0_posedge : VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SBCLKI_SBDATO1_posedge : VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SBCLKI_SBDATO2_posedge : VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SBCLKI_SBDATO3_posedge : VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SBCLKI_SBDATO4_posedge : VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SBCLKI_SBDATO5_posedge : VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SBCLKI_SBDATO6_posedge : VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SBCLKI_SBDATO7_posedge : VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SBCLKI_SBACKO_posedge : VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SBCLKI_I2CIRQ_posedge : VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SBCLKI_I2CWKUP_posedge : VitalDelayType01 := (0.000 ns, 0.000 ns);	  
------------------------added arcs--------------------------------
tpd_SCLO_SDAO_negedge: VitalDelayType01 := (0.000 ns, 0.000 ns);	
tpd_SCLO_SDAOE_negedge: VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SCLI_SDAO_negedge: VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SCLI_SDAOE_negedge: VitalDelayType01 := (0.000 ns, 0.000 ns);
------------------------------------------------------------------
----VITAL setup time
tsetup_SBRWI_SBCLKI_posedge_posedge  : VitalDelayType     := 0 ns;
tsetup_SBRWI_SBCLKI_negedge_posedge    : VitalDelayType   := 0 ns;
tsetup_SBSTBI_SBCLKI_posedge_posedge    : VitalDelayType   := 0 ns;
tsetup_SBSTBI_SBCLKI_negedge_posedge    : VitalDelayType   := 0 ns;
tsetup_SBADRI7_SBCLKI_posedge_posedge    : VitalDelayType   := 0 ns;
tsetup_SBADRI7_SBCLKI_negedge_posedge    : VitalDelayType   := 0 ns;
tsetup_SBADRI6_SBCLKI_posedge_posedge    : VitalDelayType   := 0 ns;
tsetup_SBADRI6_SBCLKI_negedge_posedge    : VitalDelayType   := 0 ns;
tsetup_SBADRI5_SBCLKI_posedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBADRI5_SBCLKI_negedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBADRI4_SBCLKI_posedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBADRI4_SBCLKI_negedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBADRI3_SBCLKI_posedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBADRI3_SBCLKI_negedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBADRI2_SBCLKI_posedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBADRI2_SBCLKI_negedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBADRI1_SBCLKI_posedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBADRI1_SBCLKI_negedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBADRI0_SBCLKI_posedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBADRI0_SBCLKI_negedge_posedge    : VitalDelayType    := 0 ns;

tsetup_SBDATI7_SBCLKI_posedge_posedge    : VitalDelayType   := 0 ns;
tsetup_SBDATI7_SBCLKI_negedge_posedge    : VitalDelayType   := 0 ns;
tsetup_SBDATI6_SBCLKI_posedge_posedge    : VitalDelayType   := 0 ns;
tsetup_SBDATI6_SBCLKI_negedge_posedge    : VitalDelayType   := 0 ns;
tsetup_SBDATI5_SBCLKI_posedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBDATI5_SBCLKI_negedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBDATI4_SBCLKI_posedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBDATI4_SBCLKI_negedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBDATI3_SBCLKI_posedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBDATI3_SBCLKI_negedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBDATI2_SBCLKI_posedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBDATI2_SBCLKI_negedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBDATI1_SBCLKI_posedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBDATI1_SBCLKI_negedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBDATI0_SBCLKI_posedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBDATI0_SBCLKI_negedge_posedge    : VitalDelayType    := 0 ns;

tsetup_SDAI_SCLO_posedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SDAI_SCLO_negedge_posedge    : VitalDelayType    := 0 ns;

tsetup_SDAI_SCLI_posedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SDAI_SCLI_negedge_posedge    : VitalDelayType    := 0 ns;


-----HOLD TIME

thold_SBRWI_SBCLKI_negedge_posedge    : VitalDelayType       := 0 ns;
thold_SBRWI_SBCLKI_posedge_posedge    : VitalDelayType        := 0 ns;
thold_SBSTBI_SBCLKI_negedge_posedge    : VitalDelayType        := 0 ns;
thold_SBSTBI_SBCLKI_posedge_posedge    : VitalDelayType        := 0 ns;
thold_SBADRI7_SBCLKI_negedge_posedge    : VitalDelayType        := 0 ns;
thold_SBADRI7_SBCLKI_posedge_posedge    : VitalDelayType        := 0 ns;
thold_SBADRI6_SBCLKI_negedge_posedge    : VitalDelayType        := 0 ns;
thold_SBADRI6_SBCLKI_posedge_posedge    : VitalDelayType        := 0 ns;
thold_SBADRI5_SBCLKI_negedge_posedge    : VitalDelayType         := 0 ns;
thold_SBADRI5_SBCLKI_posedge_posedge    : VitalDelayType         := 0 ns;
thold_SBADRI4_SBCLKI_negedge_posedge    : VitalDelayType         := 0 ns;
thold_SBADRI4_SBCLKI_posedge_posedge    : VitalDelayType         := 0 ns ;
thold_SBADRI3_SBCLKI_negedge_posedge    : VitalDelayType         := 0 ns;
thold_SBADRI3_SBCLKI_posedge_posedge    : VitalDelayType         := 0 ns;
thold_SBADRI2_SBCLKI_negedge_posedge    : VitalDelayType         := 0 ns;
thold_SBADRI2_SBCLKI_posedge_posedge    : VitalDelayType         := 0 ns;
thold_SBADRI1_SBCLKI_negedge_posedge    : VitalDelayType         := 0 ns;
thold_SBADRI1_SBCLKI_posedge_posedge    : VitalDelayType         := 0 ns;
thold_SBADRI0_SBCLKI_negedge_posedge    : VitalDelayType         := 0 ns;
thold_SBADRI0_SBCLKI_posedge_posedge    : VitalDelayType         := 0 ns;


thold_SBDATI7_SBCLKI_negedge_posedge    : VitalDelayType        := 0 ns;
thold_SBDATI7_SBCLKI_posedge_posedge    : VitalDelayType        := 0 ns;
thold_SBDATI6_SBCLKI_negedge_posedge    : VitalDelayType        := 0 ns;
thold_SBDATI6_SBCLKI_posedge_posedge    : VitalDelayType        := 0 ns;
thold_SBDATI5_SBCLKI_negedge_posedge    : VitalDelayType         := 0 ns;
thold_SBDATI5_SBCLKI_posedge_posedge    : VitalDelayType         := 0 ns;
thold_SBDATI4_SBCLKI_negedge_posedge    : VitalDelayType         := 0 ns;
thold_SBDATI4_SBCLKI_posedge_posedge    : VitalDelayType         := 0 ns ;
thold_SBDATI3_SBCLKI_negedge_posedge    : VitalDelayType         := 0 ns;
thold_SBDATI3_SBCLKI_posedge_posedge    : VitalDelayType         := 0 ns;
thold_SBDATI2_SBCLKI_negedge_posedge    : VitalDelayType         := 0 ns;
thold_SBDATI2_SBCLKI_posedge_posedge    : VitalDelayType         := 0 ns;
thold_SBDATI1_SBCLKI_negedge_posedge    : VitalDelayType         := 0 ns;
thold_SBDATI1_SBCLKI_posedge_posedge    : VitalDelayType         := 0 ns;
thold_SBDATI0_SBCLKI_negedge_posedge    : VitalDelayType         := 0 ns;
thold_SBDATI0_SBCLKI_posedge_posedge    : VitalDelayType         := 0 ns;
thold_SDAI_SCLO_posedge_posedge    : VitalDelayType    := 0 ns;
thold_SDAI_SCLO_negedge_posedge    : VitalDelayType    := 0 ns;
thold_SDAI_SCLI_posedge_posedge    : VitalDelayType    := 0 ns;
thold_SDAI_SCLI_negedge_posedge    : VitalDelayType    := 0 ns

-------SETUPHOLD WIDTH-----------
);


Port(
	    SBCLKI  : in  std_logic;
         SBRWI  : in  std_logic;
         SBSTBI  : in  std_logic;
         SBADRI7  : in  std_logic;
         SBADRI6  : in  std_logic;
         SBADRI5  : in  std_logic;
         SBADRI4  : in  std_logic;
         SBADRI3  : in  std_logic;
         SBADRI2  : in  std_logic;
         SBADRI1  : in  std_logic;
         SBADRI0  : in  std_logic;
         SBDATI7  : in  std_logic;
         SBDATI6  : in  std_logic;
         SBDATI5  : in  std_logic;
         SBDATI4  : in  std_logic;
         SBDATI3  : in  std_logic;
         SBDATI2  : in  std_logic;
         SBDATI1  : in  std_logic;
         SBDATI0  : in  std_logic;
         SCLI  : in  std_logic;
         SDAI  : in  std_logic;

        SBDATO7  : out  std_logic;
        SBDATO6  : out  std_logic;
        SBDATO5  : out  std_logic;
        SBDATO4  : out  std_logic;
        SBDATO3  : out  std_logic;
        SBDATO2  : out  std_logic;
        SBDATO1  : out  std_logic;
        SBDATO0  : out  std_logic;
        SBACKO  : out  std_logic;
        I2CIRQ  : out  std_logic;
        I2CWKUP  : out  std_logic;
        SCLO  : out  std_logic;
        SCLOE  : out  std_logic;
        SDAO  : out  std_logic;
        SDAOE  : out  std_logic
);

attribute VITAL_LEVEL0 of
    SB_I2C  : entity is true;
end SB_I2C;

architecture SB_I2C_V of SB_I2C is
  attribute VITAL_LEVEL0 of
    SB_I2C_V: architecture is true;

signal         SBCLKI_ipd  : std_ulogic := 'X';
signal         SBRWI_ipd  : std_ulogic := 'X';
signal         SBSTBI_ipd  : std_ulogic := 'X';
signal         SBADRI7_ipd  : std_ulogic := 'X';
signal         SBADRI6_ipd  : std_ulogic := 'X';
signal         SBADRI5_ipd  : std_ulogic := 'X';
signal         SBADRI4_ipd  : std_ulogic := 'X';
signal         SBADRI3_ipd  : std_ulogic := 'X';
signal         SBADRI2_ipd  : std_ulogic := 'X';
signal         SBADRI1_ipd  : std_ulogic := 'X';
signal         SBADRI0_ipd  : std_ulogic := 'X';
signal         SBDATI7_ipd  : std_ulogic := 'X';
signal         SBDATI6_ipd  : std_ulogic := 'X';
signal         SBDATI5_ipd  : std_ulogic := 'X';
signal         SBDATI4_ipd  : std_ulogic := 'X';
signal         SBDATI3_ipd  : std_ulogic := 'X';
signal         SBDATI2_ipd  : std_ulogic := 'X';
signal         SBDATI1_ipd  : std_ulogic := 'X';
signal         SBDATI0_ipd  : std_ulogic := 'X';
signal         SCLI_ipd  : std_ulogic := 'X';
signal         SDAI_ipd  : std_ulogic := 'X';
signal         SCLO_ipd  : std_ulogic := 'X';


signal        SBDATO7_sig  : std_ulogic := 'X';
signal        SBDATO6_sig  : std_ulogic := 'X';
signal        SBDATO5_sig  : std_ulogic := 'X';
signal        SBDATO4_sig  : std_ulogic := 'X';
signal        SBDATO3_sig  : std_ulogic := 'X';
signal        SBDATO2_sig  : std_ulogic := 'X';
signal        SBDATO1_sig  : std_ulogic := 'X';
signal        SBDATO0_sig  : std_ulogic := 'X';
signal        SBACKO_sig  : std_ulogic := 'X';
signal        I2CIRQ_sig  : std_ulogic := 'X';
signal        I2CWKUP_sig  : std_ulogic := 'X';
signal        SCLO_sig  : std_ulogic := 'X';
signal        SCLOE_sig  : std_ulogic := 'X';
signal        SDAO_sig  : std_ulogic := 'X';
signal        SDAOE_sig  : std_ulogic := 'X';

component SB_I2C_CORE
generic(
         I2C_SLAVE_INIT_ADDR : string := "0b1111100001";
         BUS_ADDR74 : string := "0b0001"
        );                          
port(
   SBCLKI  : in  std_logic;
         SBRWI  : in  std_logic;
         SBSTBI  : in  std_logic;
         SBADRI7  : in  std_logic;
         SBADRI6  : in  std_logic;
         SBADRI5  : in  std_logic;
         SBADRI4  : in  std_logic;
         SBADRI3  : in  std_logic;
         SBADRI2  : in  std_logic;
         SBADRI1  : in  std_logic;
         SBADRI0  : in  std_logic;
         SBDATI7  : in  std_logic;
         SBDATI6  : in  std_logic;
         SBDATI5  : in  std_logic;
         SBDATI4  : in  std_logic;
         SBDATI3  : in  std_logic;
         SBDATI2  : in  std_logic;
         SBDATI1  : in  std_logic;
         SBDATI0  : in  std_logic;
         SCLI  : in  std_logic;
         SDAI  : in  std_logic;

        SBDATO7  : out  std_logic;
        SBDATO6  : out  std_logic;
        SBDATO5  : out  std_logic;
        SBDATO4  : out  std_logic;
        SBDATO3  : out  std_logic;
        SBDATO2  : out  std_logic;
        SBDATO1  : out  std_logic;
        SBDATO0  : out  std_logic;
        SBACKO  : out  std_logic;
        I2CIRQ  : out  std_logic;
        I2CWKUP  : out  std_logic;
        SCLO  : out  std_logic;
        SCLOE  : out  std_logic;
        SDAO  : out  std_logic;
        SDAOE  : out  std_logic
);
End component;

Begin

process 
begin  
	if BUS_ADDR74 /= "0b0001" and BUS_ADDR74 /= "0b0011" then
report "ID:BUS_ADDR74: should be LLC=0b0001 or LRC=0011, otherwise there would be an error "  
severity ERROR;
end if;	 
wait ;
 end process;
	  -- SBDATO7   <= SBDATO7_zd;  
      -- SBDATO6  <= SBDATO6_zd; 
      -- SBDATO5   <= SBDATO5_zd;  
      -- SBDATO4   <= SBDATO4_zd;  
      -- SBDATO3   <= SBDATO3_zd;  
      -- SBDATO2   <= SBDATO2_zd;  
      -- SBDATO1   <= SBDATO1_zd;  
      -- SBDATO0   <= SBDATO0_zd;  
      -- SBACKO   <= SBACKO_zd;  
      -- I2CIRQ   <= I2CIRQ_zd;  
      -- I2CWKUP   <= I2CWKUP_zd;  
      SCLO   <= SCLO_sig;  
      SCLOE   <= SCLOE_sig;  
      -- SDAO   <= SDAO_zd;  
      -- SDAOE   <= SDAOE_zd;  

WireDelay : block
	Begin
VitalWireDelay	(SBCLKI_ipd,SBCLKI,tipd_SBCLKI);
VitalWireDelay	(SBRWI_ipd,SBRWI,tipd_SBRWI);
VitalWireDelay	(SBSTBI_ipd,SBSTBI,tipd_SBSTBI);
VitalWireDelay	(SBADRI7_ipd,SBADRI7,tipd_SBADRI7);
VitalWireDelay	(SBADRI6_ipd,SBADRI6,tipd_SBADRI6);
VitalWireDelay	(SBADRI5_ipd,SBADRI5,tipd_SBADRI5);
VitalWireDelay	(SBADRI4_ipd,SBADRI4,tipd_SBADRI4);
VitalWireDelay	(SBADRI3_ipd,SBADRI3,tipd_SBADRI3);
VitalWireDelay	(SBADRI2_ipd,SBADRI2,tipd_SBADRI2);
VitalWireDelay	(SBADRI1_ipd,SBADRI1,tipd_SBADRI1);
VitalWireDelay	(SBADRI0_ipd,SBADRI0,tipd_SBADRI0); 
VitalWireDelay	(SBDATI7_ipd,SBDATI7,tipd_SBDATI7);
VitalWireDelay	(SBDATI6_ipd,SBDATI6,tipd_SBDATI6);
VitalWireDelay	(SBDATI5_ipd,SBDATI5,tipd_SBDATI5);
VitalWireDelay	(SBDATI4_ipd,SBDATI4,tipd_SBDATI4);
VitalWireDelay	(SBDATI3_ipd,SBDATI3,tipd_SBDATI3);
VitalWireDelay	(SBDATI2_ipd,SBDATI2,tipd_SBDATI2);
VitalWireDelay	(SBDATI1_ipd,SBDATI1,tipd_SBDATI1);
VitalWireDelay	(SBDATI0_ipd,SBDATI0,tipd_SBDATI0);
VitalWireDelay	(SCLI_ipd,SCLI,tipd_SCLI);
VitalWireDelay	(SDAI_ipd,SDAI,tipd_SDAI);
End block;
----------------------------------------------------------------------
-- BEHAVIOR SECTION
----------------------------------------------------------------------

I2CU:SB_I2C_CORE
generic map(
            I2C_SLAVE_INIT_ADDR => I2C_SLAVE_INIT_ADDR , 
            BUS_ADDR74 => BUS_ADDR74 
            )                         
Port map(

	 SBDATO7   => SBDATO7_sig,  
      SBDATO6  => SBDATO6_sig, 
      SBDATO5   => SBDATO5_sig,  
      SBDATO4   => SBDATO4_sig,  
      SBDATO3   => SBDATO3_sig,  
      SBDATO2   => SBDATO2_sig,  
      SBDATO1   => SBDATO1_sig,  
      SBDATO0   => SBDATO0_sig,  
      SBACKO   => SBACKO_sig,  
      I2CIRQ   => I2CIRQ_sig,  
      I2CWKUP   => I2CWKUP_sig,  
      SCLO   => SCLO_sig,  
      SCLOE   => SCLOE_sig,  
      SDAO   => SDAO_sig,  
      SDAOE   => SDAOE_sig,  

	SBCLKI => SBCLKI_ipd,
	SBRWI => SBRWI_ipd,
	SBSTBI => SBSTBI_ipd,
	SBADRI7 => SBADRI7_ipd,
	SBADRI6 => SBADRI6_ipd,
	SBADRI5 => SBADRI5_ipd,
	SBADRI4 => SBADRI4_ipd,
	SBADRI3 => SBADRI3_ipd,
	SBADRI2 => SBADRI2_ipd,
	SBADRI1 => SBADRI1_ipd,
	SBADRI0 => SBADRI0_ipd,
	SBDATI7 => SBDATI7_ipd,
	SBDATI6 => SBDATI6_ipd,
	SBDATI5 => SBDATI5_ipd,
	SBDATI4 => SBDATI4_ipd,
	SBDATI3 => SBDATI3_ipd,
	SBDATI2 => SBDATI2_ipd,
	SBDATI1 => SBDATI1_ipd,
	SBDATI0 => SBDATI0_ipd,
	SCLI => SCLI_ipd,
	SDAI => SDAI_ipd
);
	
-------------------------------------------------------------------
--VITAL timing check
------------------------------------------------------------------
VITALTimingCheck : process (SBCLKI_ipd, SBRWI_ipd, SBSTBI_ipd, SBADRI7_ipd, SBADRI6_ipd, SBADRI5_ipd, SBADRI4_ipd, SBADRI3_ipd, SBADRI2_ipd, SBADRI1_ipd, SBADRI0_ipd, SBDATI7_ipd, SBDATI6_ipd, SBDATI5_ipd, SBDATI4_ipd, SBDATI3_ipd, SBDATI2_ipd, SBDATI1_ipd, SBDATI0_ipd, SCLI_ipd, SDAI_ipd)

    variable Tviol_SBRWI_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBSTBI_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SCLI_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SDATI_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBADRI7_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBADRI6_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBADRI5_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBADRI4_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBADRI3_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBADRI2_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBADRI1_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBADRI0_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBDATI7_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBDATI6_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBDATI5_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBDATI4_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBDATI3_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBDATI2_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBDATI1_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBDATI0_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SDAI_SCLO_posedge    : std_ulogic := '0';
    variable Tviol_SDAI_SCLI_posedge    : std_ulogic := '0';  
	
	
	variable Tmkr_SBRWI_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
    variable Tmkr_SBSTBI_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
	 variable Tmkr_SBRWI_SCLI_posedge     : VitalTimingDataType := VitalTimingDataInit;
    variable Tmkr_SDATI_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
    variable Tmkr_SBADRI7_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
    variable Tmkr_SBADRI6_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
    variable Tmkr_SBADRI5_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
	 variable Tmkr_SBADRI4_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
    variable Tmkr_SBADRI3_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
    variable Tmkr_SBADRI2_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
    variable Tmkr_SBADRI1_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
    variable Tmkr_SBADRI0_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
	 variable Tmkr_SBDATI7_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
    variable Tmkr_SBDATI6_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
    variable Tmkr_SBDATI5_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
	 variable Tmkr_SBDATI4_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
    variable Tmkr_SBDATI3_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
    variable Tmkr_SBDATI2_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
    variable Tmkr_SBDATI1_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
    variable Tmkr_SBDATI0_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_SDAI_SCLO_posedge     : VitalTimingDataType := VitalTimingDataInit;
    variable Tmkr_SDAI_SCLI_posedge     : VitalTimingDataType := VitalTimingDataInit; 


begin
if (TimingChecksOn) then
      VitalSetupHoldCheck (
        Violation      => Tviol_SBRWI_SBCLKI_posedge,
        TimingData     => Tmkr_SBRWI_SBCLKI_posedge,
        TestSignal     => SBRWI_ipd,
        TestSignalName => "SBRWI",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBRWI_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBRWI_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBRWI_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBRWI_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);
 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBSTBI_SBCLKI_posedge,
        TimingData     => Tmkr_SBSTBI_SBCLKI_posedge,
        TestSignal     => SBSTBI_ipd,
        TestSignalName => "SBSTBI",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBSTBI_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBSTBI_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBSTBI_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBSTBI_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);
 		 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBADRI7_SBCLKI_posedge,
        TimingData     => Tmkr_SBADRI7_SBCLKI_posedge,
        TestSignal     => SBADRI7_ipd,
        TestSignalName => "SBADRI7",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBADRI7_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBADRI7_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBADRI7_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBADRI7_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);		
 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBADRI6_SBCLKI_posedge,
        TimingData     => Tmkr_SBADRI6_SBCLKI_posedge,
        TestSignal     => SBADRI6_ipd,
        TestSignalName => "SBADRI6",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBADRI6_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBADRI6_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBADRI6_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBADRI6_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);		

		 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBADRI5_SBCLKI_posedge,
        TimingData     => Tmkr_SBADRI5_SBCLKI_posedge,
        TestSignal     => SBADRI5_ipd,
        TestSignalName => "SBADRI5",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBADRI5_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBADRI5_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBADRI5_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBADRI5_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);		
		
 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBADRI4_SBCLKI_posedge,
        TimingData     => Tmkr_SBADRI4_SBCLKI_posedge,
        TestSignal     => SBADRI4_ipd,
        TestSignalName => "SBADRI4",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBADRI4_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBADRI4_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBADRI4_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBADRI4_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);	
 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBADRI3_SBCLKI_posedge,
        TimingData     => Tmkr_SBADRI3_SBCLKI_posedge,
        TestSignal     => SBADRI3_ipd,
        TestSignalName => "SBADRI3",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBADRI3_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBADRI3_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBADRI3_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBADRI3_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);		
 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBADRI2_SBCLKI_posedge,
        TimingData     => Tmkr_SBADRI2_SBCLKI_posedge,
        TestSignal     => SBADRI2_ipd,
        TestSignalName => "SBADRI2",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBADRI2_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBADRI2_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBADRI2_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBADRI2_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);
 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBADRI1_SBCLKI_posedge,
        TimingData     => Tmkr_SBADRI1_SBCLKI_posedge,
        TestSignal     => SBADRI1_ipd,
        TestSignalName => "SBADRI1",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBADRI1_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBADRI1_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBADRI1_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBADRI1_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);	
 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBADRI0_SBCLKI_posedge,
        TimingData     => Tmkr_SBADRI0_SBCLKI_posedge,
        TestSignal     => SBADRI0_ipd,
        TestSignalName => "SBADRI0",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBADRI0_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBADRI0_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBADRI0_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBADRI0_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);		
		 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBDATI7_SBCLKI_posedge,
        TimingData     => Tmkr_SBDATI7_SBCLKI_posedge,
        TestSignal     => SBDATI7_ipd,
        TestSignalName => "SBDATI7",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBDATI7_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBDATI7_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBDATI7_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBDATI7_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);		
 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBDATI6_SBCLKI_posedge,
        TimingData     => Tmkr_SBDATI6_SBCLKI_posedge,
        TestSignal     => SBDATI6_ipd,
        TestSignalName => "SBDATI6",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBDATI6_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBDATI6_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBDATI6_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBDATI6_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);		

		 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBDATI5_SBCLKI_posedge,
        TimingData     => Tmkr_SBDATI5_SBCLKI_posedge,
        TestSignal     => SBDATI5_ipd,
        TestSignalName => "SBDATI5",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBDATI5_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBDATI5_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBDATI5_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBDATI5_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);		
		
 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBDATI4_SBCLKI_posedge,
        TimingData     => Tmkr_SBDATI4_SBCLKI_posedge,
        TestSignal     => SBDATI4_ipd,
        TestSignalName => "SBDATI4",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBDATI4_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBDATI4_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBDATI4_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBDATI4_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);	
 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBDATI3_SBCLKI_posedge,
        TimingData     => Tmkr_SBDATI3_SBCLKI_posedge,
        TestSignal     => SBDATI3_ipd,
        TestSignalName => "SBDATI3",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBDATI3_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBDATI3_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBDATI3_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBDATI3_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);		
 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBDATI2_SBCLKI_posedge,
        TimingData     => Tmkr_SBDATI2_SBCLKI_posedge,
        TestSignal     => SBDATI2_ipd,
        TestSignalName => "SBDATI2",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBDATI2_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBDATI2_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBDATI2_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBDATI2_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);
 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBDATI1_SBCLKI_posedge,
        TimingData     => Tmkr_SBDATI1_SBCLKI_posedge,
        TestSignal     => SBDATI1_ipd,
        TestSignalName => "SBDATI1",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBDATI1_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBDATI1_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBDATI1_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBDATI1_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);	
 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBDATI0_SBCLKI_posedge,
        TimingData     => Tmkr_SBDATI0_SBCLKI_posedge,
        TestSignal     => SBDATI0_ipd,
        TestSignalName => "SBDATI0",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBDATI0_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBDATI0_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBDATI0_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBDATI0_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);	
	VitalSetupHoldCheck (
        Violation      => Tviol_SDAI_SCLO_posedge,
        TimingData     => Tmkr_SDAI_SCLO_posedge,
        TestSignal     => SDAI_ipd,
        TestSignalName => "SDAI",
        RefSignal      => SCLO_ipd,
        RefSignalName  => "SCLO",
        SetupHigh      => tsetup_SDAI_SCLO_posedge_posedge,
        SetupLow       => tsetup_SDAI_SCLO_negedge_posedge,
        HoldLow        => thold_SDAI_SCLO_negedge_posedge,
        HoldHigh       => thold_SDAI_SCLO_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);			
		
	VitalSetupHoldCheck (
        Violation      => Tviol_SDAI_SCLI_posedge,
        TimingData     => Tmkr_SDAI_SCLI_posedge,
        TestSignal     => SDAI_ipd,
        TestSignalName => "SDAI",
        RefSignal      => SCLI_ipd,
        RefSignalName  => "SCLI",
        SetupHigh      => tsetup_SDAI_SCLI_posedge_posedge,
        SetupLow       => tsetup_SDAI_SCLI_negedge_posedge,
        HoldLow        => thold_SDAI_SCLI_negedge_posedge,
        HoldHigh       => thold_SDAI_SCLI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);		


end if;
end process;

VITALPathDelay   : process (SBCLKI_ipd, SBRWI_ipd, SBSTBI_ipd, SCLI_ipd, 
SDAI_ipd,SBDATO7_sig,SBDATO6_sig,SBDATO5_sig, SBDATO4_sig,SBDATO3_sig,SBDATO2_sig,SBDATO1_sig, SBDATO0_sig,SBACKO_sig,I2CIRQ_sig,I2CWKUP_sig,SCLO_sig,  
SDAO_sig,SDAOE_sig)
variable SBDATO7_GlitchData : VitalGlitchDataType;  
variable SBDATO6_GlitchData : VitalGlitchDataType;
variable SBDATO5_GlitchData : VitalGlitchDataType;
variable SBDATO4_GlitchData : VitalGlitchDataType;
variable SBDATO3_GlitchData : VitalGlitchDataType;
variable SBDATO2_GlitchData : VitalGlitchDataType;
variable SBDATO1_GlitchData : VitalGlitchDataType;
variable SBDATO0_GlitchData : VitalGlitchDataType;
variable SBACKO_GlitchData : VitalGlitchDataType;
variable I2CIRQ_GlitchData : VitalGlitchDataType;
variable I2CWKUP_GlitchData : VitalGlitchDataType;
variable SCLO_GlitchData : VitalGlitchDataType;
variable SCLOE_GlitchData : VitalGlitchDataType;
variable SDAO_GlitchData : VitalGlitchDataType;
variable SDAOE_GlitchData : VitalGlitchDataType;
		 
variable        SBDATO7_zd  : std_ulogic := 'X';
variable        SBDATO6_zd  : std_ulogic := 'X';
variable        SBDATO5_zd  : std_ulogic := 'X';
variable        SBDATO4_zd  : std_ulogic := 'X';
variable        SBDATO3_zd  : std_ulogic := 'X';
variable        SBDATO2_zd  : std_ulogic := 'X';
variable        SBDATO1_zd  : std_ulogic := 'X';
variable        SBDATO0_zd  : std_ulogic := 'X';
variable        SBACKO_zd  : std_ulogic := 'X';
variable        I2CIRQ_zd  : std_ulogic := 'X';
variable        I2CWKUP_zd  : std_ulogic := 'X';
variable        SCLO_zd  : std_ulogic := 'X';
variable        SCLOE_zd  : std_ulogic := 'X';
variable        SDAO_zd  : std_ulogic := 'X';
variable        SDAOE_zd  : std_ulogic := 'X';

begin	  
	
	SDAO_zd := SDAO_sig;	
	        SBDATO7_zd  := SBDATO7_sig;
        SBDATO6_zd  := SBDATO6_sig;
        SBDATO5_zd  := SBDATO5_sig;
        SBDATO4_zd  := SBDATO4_sig;
        SBDATO3_zd  := SBDATO3_sig;
        SBDATO2_zd  := SBDATO2_sig;
        SBDATO1_zd  := SBDATO1_sig;
        SBDATO0_zd  := SBDATO0_sig;
        SBACKO_zd  := SBACKO_sig;
        I2CIRQ_zd  := I2CIRQ_sig;
        I2CWKUP_zd  := I2CWKUP_sig;
        SCLO_zd  := SCLO_sig;
        SCLOE_zd  := SCLOE_sig;
        SDAO_zd  := SDAO_sig;
        SDAOE_zd  := SDAOE_sig;
	
  VitalPathDelay01 (
      OutSignal                 => SBDATO7,
      GlitchData                => SBDATO7_GlitchData,
      OutSignalName             => "SBDATO7",
      OutTemp                   => SBDATO7_zd,
      Paths                     => (0 => (SBCLKI_ipd'last_event, tpd_SBCLKI_SBDATO7_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);	 
VitalPathDelay01 (
      OutSignal                 => SBDATO6,
      GlitchData                => SBDATO6_GlitchData,
      OutSignalName             => "SBDATO6",
      OutTemp                   => SBDATO6_zd,
      Paths                     => (0 => (SBCLKI_ipd'last_event, tpd_SBCLKI_SBDATO6_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

  VitalPathDelay01 (
      OutSignal                 => SBDATO5,
      GlitchData                => SBDATO5_GlitchData,
      OutSignalName             => "SBDATO5",
      OutTemp                   => SBDATO5_zd,
      Paths                     => (0 => (SBCLKI_ipd'last_event, tpd_SBCLKI_SBDATO5_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

  VitalPathDelay01 (
      OutSignal                 => SBDATO4,
      GlitchData                => SBDATO4_GlitchData,
      OutSignalName             => "SBDATO4",
      OutTemp                   => SBDATO4_zd,
      Paths                     => (0 => (SBCLKI_ipd'last_event, tpd_SBCLKI_SBDATO4_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

  VitalPathDelay01 (
      OutSignal                 => SBDATO3,
      GlitchData                => SBDATO3_GlitchData,
      OutSignalName             => "SBDATO3",
      OutTemp                   => SBDATO3_zd,
      Paths                     => (0 => (SBCLKI_ipd'last_event, tpd_SBCLKI_SBDATO3_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);


  VitalPathDelay01 (
      OutSignal                 => SBDATO2,
      GlitchData                => SBDATO2_GlitchData,
      OutSignalName             => "SBDATO2",
      OutTemp                   => SBDATO2_zd,
      Paths                     => (0 => (SBCLKI_ipd'last_event, tpd_SBCLKI_SBDATO2_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

  VitalPathDelay01 (
      OutSignal                 => SBDATO1,
      GlitchData                => SBDATO1_GlitchData,
      OutSignalName             => "SBDATO1",
      OutTemp                   => SBDATO1_zd,
      Paths                     => (0 => (SBCLKI_ipd'last_event, tpd_SBCLKI_SBDATO1_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

  VitalPathDelay01 (
      OutSignal                 => SBDATO0,
      GlitchData                => SBDATO0_GlitchData,
      OutSignalName             => "SBDATO0",
      OutTemp                   => SBDATO0_zd,
      Paths                     => (0 => (SBCLKI_ipd'last_event, tpd_SBCLKI_SBDATO0_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

  VitalPathDelay01 (
      OutSignal                 => SBACKO,
      GlitchData                => SBACKO_GlitchData,
      OutSignalName             => "SBACKO",
      OutTemp                   => SBACKO_zd,
      Paths                     => (0 => (SBCLKI_ipd'last_event, tpd_SBCLKI_SBACKO_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

VitalPathDelay01 (
      OutSignal                 => I2CIRQ,
      GlitchData                => I2CIRQ_GlitchData,
      OutSignalName             => "I2CIRQ",
      OutTemp                   => I2CIRQ_zd,
      Paths                     => (0 => (SBCLKI_ipd'last_event, tpd_SBCLKI_I2CIRQ_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

VitalPathDelay01 (
      OutSignal                 => I2CWKUP,
      GlitchData                => I2CWKUP_GlitchData,
      OutSignalName             => "I2CWKUP",
      OutTemp                   => I2CWKUP_zd,
      Paths                     => (0 => (SBCLKI_ipd'last_event, tpd_SBCLKI_I2CWKUP_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);


VitalPathDelay01 (
      OutSignal                 => SDAOE,
      GlitchData                => SDAOE_GlitchData,
      OutSignalName             => "SDAOE",
      OutTemp                   => SDAOE_zd,
      Paths                     => (0 => (SCLO_ipd'last_event, tpd_SCLO_SDAOE_negedge, true),
	 								1 => (SCLI_ipd'last_event, tpd_SCLI_SDAOE_negedge, true),
	  								2 => (SCLO_ipd'last_event, tpd_SCLO_SDAOE_posedge, true),
	  								3 => (SCLI_ipd'last_event, tpd_SCLI_SDAOE_posedge, true)),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

VitalPathDelay01 (
      OutSignal                 => SDAO,
      GlitchData                => SDAO_GlitchData,
      OutSignalName             => "SDAO",
      OutTemp                   => SDAO_zd,
      Paths                     => (0 => (SCLI_ipd'last_event, tpd_SCLI_SDAO_negedge, true),	
	  								1 => (SCLO_ipd'last_event, tpd_SCLI_SDAO_posedge, true),
	  								2 => (SCLO_ipd'last_event, tpd_SCLO_SDAO_posedge, true),
									3 => (SCLO_ipd'last_event, tpd_SCLO_SDAO_negedge, true)
									),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);



  end process VITALPathDelay;

end SB_I2C_V;

-----------------------------------------------
----       SB_SPI 			------
----------------------------------------------
library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use IEEE.Vital_Primitives.all;
use IEEE.VITAL_Timing.all;
library WORK;
use WORK.vcomponent_vital.all;

entity  SB_SPI  is 
--define kinds of delay timing paras default value
	generic(
	BUS_ADDR74 : string := "0b0000" ;
	---------------------------------------------------------------
----VITAL PARAMETER	
--	------------------------------------------
TimingChecksOn  : boolean := true;
	Xon   : boolean := true;			    
    	MsgOn : boolean := false;
	--Vital path delay
Tipd_SBCLKI : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBRWI : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBSTBI : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBADRI7 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBADRI6 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBADRI5 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBADRI4 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBADRI3 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBADRI2 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBADRI1 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBADRI0 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBDATI7 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBDATI6 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBDATI5 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBDATI4 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBDATI3 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBDATI2 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBDATI1 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SBDATI0 : VitalDelayType01 := (0 ns, 0 ns);
Tipd_MI : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SI : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SCKI : VitalDelayType01 := (0 ns, 0 ns);
Tipd_SCSNI : VitalDelayType01 := (0 ns, 0 ns);

--Vital path delay
tpd_SCKO_MO_posedge : VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SCKO_MO_negedge : VitalDelayType01 := (0.000 ns, 0.000 ns);	-----------------
tpd_SCKO_MOE_posedge : VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SCKO_MCSNO3_posedge : VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SCKO_MCSNO2_posedge: VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SCKO_MCSNO1_posedge: VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SCKO_MCSNO0_posedge: VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SCKO_MCSNOE3_posedge: VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SCKO_MCSNOE2_posedge: VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SCKO_MCSNOE1_posedge: VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SCKO_MCSNOE0_posedge: VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SCKI_SO_posedge: VitalDelayType01 := (0.000 ns, 0.000 ns);	
tpd_SCKI_SO_negedge: VitalDelayType01 := (0.000 ns, 0.000 ns); ----------------
tpd_SCKI_SOE_posedge: VitalDelayType01 := (0.000 ns, 0.000 ns);
--Vital clk-to-output path delay
--tpd_SBCLKI_SCKO : VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SBCLKI_SBDATO0_posedge : VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SBCLKI_SBDATO1_posedge : VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SBCLKI_SBDATO2_posedge : VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SBCLKI_SBDATO3_posedge : VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SBCLKI_SBDATO4_posedge : VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SBCLKI_SBDATO5_posedge : VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SBCLKI_SBDATO6_posedge : VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SBCLKI_SBDATO7_posedge : VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SBCLKI_SBACKO_posedge : VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SBCLKI_SPIIRQ_posedge : VitalDelayType01 := (0.000 ns, 0.000 ns);
tpd_SBCLKI_SPIWKUP_posedge : VitalDelayType01 := (0.000 ns, 0.000 ns); 

----VITAL setup time
tsetup_SBRWI_SBCLKI_posedge_posedge  : VitalDelayType     := 0 ns;
tsetup_SBRWI_SBCLKI_negedge_posedge    : VitalDelayType   := 0 ns;
tsetup_SBSTBI_SBCLKI_posedge_posedge    : VitalDelayType   := 0 ns;
tsetup_SBSTBI_SBCLKI_negedge_posedge    : VitalDelayType   := 0 ns;
tsetup_SBADRI7_SBCLKI_posedge_posedge    : VitalDelayType   := 0 ns;
tsetup_SBADRI7_SBCLKI_negedge_posedge    : VitalDelayType   := 0 ns;
tsetup_SBADRI6_SBCLKI_posedge_posedge    : VitalDelayType   := 0 ns;
tsetup_SBADRI6_SBCLKI_negedge_posedge    : VitalDelayType   := 0 ns;
tsetup_SBADRI5_SBCLKI_posedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBADRI5_SBCLKI_negedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBADRI4_SBCLKI_posedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBADRI4_SBCLKI_negedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBADRI3_SBCLKI_posedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBADRI3_SBCLKI_negedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBADRI2_SBCLKI_posedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBADRI2_SBCLKI_negedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBADRI1_SBCLKI_posedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBADRI1_SBCLKI_negedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBADRI0_SBCLKI_posedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBADRI0_SBCLKI_negedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBDATI7_SBCLKI_posedge_posedge    : VitalDelayType   := 0 ns;
tsetup_SBDATI7_SBCLKI_negedge_posedge    : VitalDelayType   := 0 ns;
tsetup_SBDATI6_SBCLKI_posedge_posedge    : VitalDelayType   := 0 ns;
tsetup_SBDATI6_SBCLKI_negedge_posedge    : VitalDelayType   := 0 ns;
tsetup_SBDATI5_SBCLKI_posedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBDATI5_SBCLKI_negedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBDATI4_SBCLKI_posedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBDATI4_SBCLKI_negedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBDATI3_SBCLKI_posedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBDATI3_SBCLKI_negedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBDATI2_SBCLKI_posedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBDATI2_SBCLKI_negedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBDATI1_SBCLKI_posedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBDATI1_SBCLKI_negedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBDATI0_SBCLKI_posedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SBDATI0_SBCLKI_negedge_posedge    : VitalDelayType    := 0 ns;
tsetup_MI_SCKO_posedge_posedge    : VitalDelayType    := 0 ns;
tsetup_MI_SCKO_negedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SI_SCKI_posedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SI_SCKI_negedge_posedge    : VitalDelayType    := 0 ns;								 
tsetup_SCSNI_SCKI_posedge_posedge    : VitalDelayType    := 0 ns;
tsetup_SCSNI_SCKI_negedge_posedge    : VitalDelayType    := 0 ns; 
---------------------------added---------------------------------
tsetup_MI_SCKO_posedge_negedge    : VitalDelayType    := 0 ns;
tsetup_MI_SCKO_negedge_negedge    : VitalDelayType    := 0 ns;
tsetup_SI_SCKI_posedge_negedge    : VitalDelayType    := 0 ns;
tsetup_SI_SCKI_negedge_negedge    : VitalDelayType    := 0 ns;								 
tsetup_SCSNI_SCKI_posedge_negedge    : VitalDelayType    := 0 ns;
tsetup_SCSNI_SCKI_negedge_negedge    : VitalDelayType    := 0 ns; 
-----------------------------------------------------------------

-----HOLD TIME

thold_SBRWI_SBCLKI_negedge_posedge    : VitalDelayType       := 0 ns;
thold_SBRWI_SBCLKI_posedge_posedge    : VitalDelayType        := 0 ns;
thold_SBSTBI_SBCLKI_negedge_posedge    : VitalDelayType        := 0 ns;
thold_SBSTBI_SBCLKI_posedge_posedge    : VitalDelayType        := 0 ns;
thold_SBADRI7_SBCLKI_negedge_posedge    : VitalDelayType        := 0 ns;
thold_SBADRI7_SBCLKI_posedge_posedge    : VitalDelayType        := 0 ns;
thold_SBADRI6_SBCLKI_negedge_posedge    : VitalDelayType        := 0 ns;
thold_SBADRI6_SBCLKI_posedge_posedge    : VitalDelayType        := 0 ns;
thold_SBADRI5_SBCLKI_negedge_posedge    : VitalDelayType         := 0 ns;
thold_SBADRI5_SBCLKI_posedge_posedge    : VitalDelayType         := 0 ns;
thold_SBADRI4_SBCLKI_negedge_posedge    : VitalDelayType         := 0 ns;
thold_SBADRI4_SBCLKI_posedge_posedge    : VitalDelayType         := 0 ns ;
thold_SBADRI3_SBCLKI_negedge_posedge    : VitalDelayType         := 0 ns;
thold_SBADRI3_SBCLKI_posedge_posedge    : VitalDelayType         := 0 ns;
thold_SBADRI2_SBCLKI_negedge_posedge    : VitalDelayType         := 0 ns;
thold_SBADRI2_SBCLKI_posedge_posedge    : VitalDelayType         := 0 ns;
thold_SBADRI1_SBCLKI_negedge_posedge    : VitalDelayType         := 0 ns;
thold_SBADRI1_SBCLKI_posedge_posedge    : VitalDelayType         := 0 ns;
thold_SBADRI0_SBCLKI_negedge_posedge    : VitalDelayType         := 0 ns;
thold_SBADRI0_SBCLKI_posedge_posedge    : VitalDelayType         := 0 ns;


thold_SBDATI7_SBCLKI_negedge_posedge    : VitalDelayType        := 0 ns;
thold_SBDATI7_SBCLKI_posedge_posedge    : VitalDelayType        := 0 ns;
thold_SBDATI6_SBCLKI_negedge_posedge    : VitalDelayType        := 0 ns;
thold_SBDATI6_SBCLKI_posedge_posedge    : VitalDelayType        := 0 ns;
thold_SBDATI5_SBCLKI_negedge_posedge    : VitalDelayType         := 0 ns;
thold_SBDATI5_SBCLKI_posedge_posedge    : VitalDelayType         := 0 ns;
thold_SBDATI4_SBCLKI_negedge_posedge    : VitalDelayType         := 0 ns;
thold_SBDATI4_SBCLKI_posedge_posedge    : VitalDelayType         := 0 ns ;
thold_SBDATI3_SBCLKI_negedge_posedge    : VitalDelayType         := 0 ns;
thold_SBDATI3_SBCLKI_posedge_posedge    : VitalDelayType         := 0 ns;
thold_SBDATI2_SBCLKI_negedge_posedge    : VitalDelayType         := 0 ns;
thold_SBDATI2_SBCLKI_posedge_posedge    : VitalDelayType         := 0 ns;
thold_SBDATI1_SBCLKI_negedge_posedge    : VitalDelayType         := 0 ns;
thold_SBDATI1_SBCLKI_posedge_posedge    : VitalDelayType         := 0 ns;
thold_SBDATI0_SBCLKI_negedge_posedge    : VitalDelayType         := 0 ns;
thold_SBDATI0_SBCLKI_posedge_posedge    : VitalDelayType         := 0 ns;
thold_MI_SCKO_posedge_posedge    : VitalDelayType    := 0 ns;
thold_MI_SCKO_negedge_posedge    : VitalDelayType    := 0 ns;					  
thold_SI_SCKI_posedge_posedge    : VitalDelayType    := 0 ns;
thold_SI_SCKI_negedge_posedge    : VitalDelayType    := 0 ns;
thold_SCSNI_SCKI_posedge_posedge    : VitalDelayType    := 0 ns;
thold_SCSNI_SCKI_negedge_posedge    : VitalDelayType    := 0 ns;
---------------------------added---------------------------------
thold_MI_SCKO_posedge_negedge    : VitalDelayType    := 0 ns;
thold_MI_SCKO_negedge_negedge    : VitalDelayType    := 0 ns;
thold_SI_SCKI_posedge_negedge    : VitalDelayType    := 0 ns;
thold_SI_SCKI_negedge_negedge    : VitalDelayType    := 0 ns;								 
thold_SCSNI_SCKI_posedge_negedge    : VitalDelayType    := 0 ns;
thold_SCSNI_SCKI_negedge_negedge    : VitalDelayType    := 0 ns 
-----------------------------------------------------------------
--
-------SETUPHOLD WIDTH-----------
);


Port(
	    SBCLKI  : in  std_logic;
         SBRWI  : in  std_logic;
         SBSTBI  : in  std_logic;
         SBADRI7  : in  std_logic;
         SBADRI6  : in  std_logic;
         SBADRI5  : in  std_logic;
         SBADRI4  : in  std_logic;
         SBADRI3  : in  std_logic;
         SBADRI2  : in  std_logic;
         SBADRI1  : in  std_logic;
         SBADRI0  : in  std_logic;
         SBDATI7  : in  std_logic;
         SBDATI6  : in  std_logic;
         SBDATI5  : in  std_logic;
         SBDATI4  : in  std_logic;
         SBDATI3  : in  std_logic;
         SBDATI2  : in  std_logic;
         SBDATI1  : in  std_logic;
         SBDATI0  : in  std_logic;
         MI  : in  std_logic;
         SI  : in  std_logic;
	      SCKI: in  std_logic;
         SCSNI : in  std_logic;


        SBDATO7  : out  std_logic;
        SBDATO6  : out  std_logic;
        SBDATO5  : out  std_logic;
        SBDATO4  : out  std_logic;
        SBDATO3  : out  std_logic;
        SBDATO2  : out  std_logic;
        SBDATO1  : out  std_logic;
        SBDATO0  : out  std_logic;
        SBACKO  : out  std_logic;
        SPIIRQ  : out  std_logic;
        SPIWKUP  : out  std_logic;
        SO  : out  std_logic;
        SOE  : out  std_logic;
        MO  : out  std_logic;
        MOE  : out  std_logic;
        SCKO  : out  std_logic;
        SCKOE  : out  std_logic;
        MCSNO3  : out  std_logic;
       
		MCSNO2  : out  std_logic;
		MCSNO1  : out  std_logic;
		MCSNO0  : out  std_logic;
		MCSNOE3  : out  std_logic;
		MCSNOE2  : out  std_logic;
		MCSNOE1  : out  std_logic;
		MCSNOE0  : out  std_logic


);

attribute VITAL_LEVEL0 of
   SB_SPI  : entity is true;
end SB_SPI;

architecture SB_SPI_V of SB_SPI is
  attribute VITAL_LEVEL0 of
    SB_SPI_V: architecture is true;

component SB_SPI_CORE
  generic(
                  BUS_ADDR74 : string := "0b0000"
         ); 
port(
   SBCLKI  : in  std_logic;
         SBRWI  : in  std_logic;
         SBSTBI  : in  std_logic;
         SBADRI7  : in  std_logic;
         SBADRI6  : in  std_logic;
         SBADRI5  : in  std_logic;
         SBADRI4  : in  std_logic;
         SBADRI3  : in  std_logic;
         SBADRI2  : in  std_logic;
         SBADRI1  : in  std_logic;
         SBADRI0  : in  std_logic;
         SBDATI7  : in  std_logic;
         SBDATI6  : in  std_logic;
         SBDATI5  : in  std_logic;
         SBDATI4  : in  std_logic;
         SBDATI3  : in  std_logic;
         SBDATI2  : in  std_logic;
         SBDATI1  : in  std_logic;
         SBDATI0  : in  std_logic;
         MI  : in  std_logic;
         SI  : in  std_logic;
		 SCKI  : in  std_logic;
         SCSNI : in  std_logic;
	

        SBDATO7  : out  std_logic;
        SBDATO6  : out  std_logic;
        SBDATO5  : out  std_logic;
        SBDATO4  : out  std_logic;
        SBDATO3  : out  std_logic;
        SBDATO2  : out  std_logic;
        SBDATO1  : out  std_logic;
        SBDATO0  : out  std_logic;
        SBACKO  : out  std_logic;
        SPIIRQ  : out  std_logic;
        SPIWKUP  : out  std_logic;
        SO  : out  std_logic;
        SOE  : out  std_logic;
        MO  : out  std_logic;
        MOE  : out  std_logic;
        SCKO  : out  std_logic;
        SCKOE  : out  std_logic;
        MCSNO3  : out  std_logic;
        MCSNO2  : out  std_logic;
        MCSNO1  : out  std_logic;
        MCSNO0  : out  std_logic;
        MCSNOE3  : out  std_logic;
        MCSNOE2  : out  std_logic;
	     MCSNOE1 : out  std_logic;
        MCSNOE0  : out  std_logic

);
End component;

signal         SBCLKI_ipd  : std_ulogic := 'X';
signal         SBRWI_ipd  : std_ulogic := 'X';
signal         SBSTBI_ipd  : std_ulogic := 'X';
signal         SBADRI7_ipd  : std_ulogic := 'X';
signal         SBADRI6_ipd  : std_ulogic := 'X';
signal         SBADRI5_ipd  : std_ulogic := 'X';
signal         SBADRI4_ipd  : std_ulogic := 'X';
signal         SBADRI3_ipd  : std_ulogic := 'X';
signal         SBADRI2_ipd  : std_ulogic := 'X';
signal         SBADRI1_ipd  : std_ulogic := 'X';
signal         SBADRI0_ipd  : std_ulogic := 'X';
signal         SBDATI7_ipd  : std_ulogic := 'X';
signal         SBDATI6_ipd  : std_ulogic := 'X';
signal         SBDATI5_ipd  : std_ulogic := 'X';
signal         SBDATI4_ipd  : std_ulogic := 'X';
signal         SBDATI3_ipd  : std_ulogic := 'X';
signal         SBDATI2_ipd  : std_ulogic := 'X';
signal         SBDATI1_ipd  : std_ulogic := 'X';
signal         SBDATI0_ipd  : std_ulogic := 'X';
signal         MI_ipd  : std_ulogic := 'X';
signal         SI_ipd  : std_ulogic := 'X';
signal         SCKI_ipd  : std_ulogic := 'X';
signal         SCSNI_ipd  : std_ulogic := 'X'; 					 

--signal         SCKO_zd  : std_ulogic := 'X';
signal        SBDATO7_zd  : std_ulogic := 'X';
signal        SBDATO6_zd  : std_ulogic := 'X';
signal        SBDATO5_zd  : std_ulogic := 'X';
signal        SBDATO4_zd  : std_ulogic := 'X';
signal        SBDATO3_zd  : std_ulogic := 'X';
signal        SBDATO2_zd  : std_ulogic := 'X';
signal        SBDATO1_zd  : std_ulogic := 'X';
signal        SBDATO0_zd  : std_ulogic := 'X';
signal        SBACKO_zd  : std_ulogic := 'X';
signal        SPIIRQ_zd  : std_ulogic := 'X';
signal        SPIWKUP_zd  : std_ulogic := 'X';
signal        SO_zd  : std_ulogic := 'X';
signal        SOE_zd  : std_ulogic := 'X';
signal        MO_zd  : std_ulogic := 'X';
signal        MOE_zd  : std_ulogic := 'X';
signal        SCKO_zd  : std_ulogic := 'X';
signal        SCKOE_zd  : std_ulogic := 'X';
signal        MCSNO3_zd  : std_ulogic := 'X';
signal        MCSNO2_zd  : std_ulogic := 'X';
signal        MCSNO1_zd  : std_ulogic := 'X';
signal        MCSNO0_zd  : std_ulogic := 'X';
signal        MCSNOE3_zd  : std_ulogic := 'X';
signal        MCSNOE2_zd  : std_ulogic := 'X';
signal        MCSNOE1_zd  : std_ulogic := 'X';
signal        MCSNOE0_zd  : std_ulogic := 'X';

begin  
			   -- SBDATO7  <=SBDATO7_zd;
               -- SBDATO6  <=SBDATO6_zd;
               -- SBDATO5  <=SBDATO5_zd;	
               -- SBDATO4  <=SBDATO4_zd;
               -- SBDATO3  <=SBDATO3_zd;
               -- SBDATO2  <=SBDATO2_zd;
               -- SBDATO1  <=SBDATO1_zd;
               -- SBDATO0  <=SBDATO0_zd;
               -- SBACKO  <=SBACKO_zd;
               -- SPIIRQ  <=SPIIRQ_zd;
               -- SPIWKUP  <=SPIWKUP_zd;
               -- SO  <=SO_zd;
               -- SOE  <=SOE_zd;
               -- MO  <=MO_zd;
               -- MOE  <=MOE_zd;
               SCKO  <=SCKO_zd;
               SCKOE  <=SCKOE_zd;
               -- MCSNO3  <=MCSNO3_zd;
               -- MCSNO2  <=MCSNO2_zd;
               -- MCSNO1  <=MCSNO1_zd;
               -- MCSNO0  <=MCSNO0_zd;
               -- MCSNOE3  <=MCSNOE3_zd;
               -- MCSNOE2  <=MCSNOE2_zd;
               -- MCSNOE1  <=MCSNOE1_zd;
               -- MCSNOE0  <=MCSNOE0_zd;	
WireDelay : block
	Begin
VitalWireDelay	(SBCLKI_ipd,SBCLKI,tipd_SBCLKI);
VitalWireDelay	(SBRWI_ipd,SBRWI,tipd_SBRWI);
VitalWireDelay	(SBSTBI_ipd,SBSTBI,tipd_SBSTBI);
VitalWireDelay	(SBADRI7_ipd,SBADRI7,tipd_SBADRI7);
VitalWireDelay	(SBADRI6_ipd,SBADRI6,tipd_SBADRI6);
VitalWireDelay	(SBADRI5_ipd,SBADRI5,tipd_SBADRI5);
VitalWireDelay	(SBADRI4_ipd,SBADRI4,tipd_SBADRI4);
VitalWireDelay	(SBADRI3_ipd,SBADRI3,tipd_SBADRI3);
VitalWireDelay	(SBADRI2_ipd,SBADRI2,tipd_SBADRI2);
VitalWireDelay	(SBADRI1_ipd,SBADRI1,tipd_SBADRI1);
VitalWireDelay	(SBADRI0_ipd,SBADRI0,tipd_SBADRI0); 
VitalWireDelay	(SBDATI7_ipd,SBDATI7,tipd_SBDATI7);
VitalWireDelay	(SBDATI6_ipd,SBDATI6,tipd_SBDATI6);
VitalWireDelay	(SBDATI5_ipd,SBDATI5,tipd_SBDATI5);
VitalWireDelay	(SBDATI4_ipd,SBDATI4,tipd_SBDATI4);
VitalWireDelay	(SBDATI3_ipd,SBDATI3,tipd_SBDATI3);
VitalWireDelay	(SBDATI2_ipd,SBDATI2,tipd_SBDATI2);
VitalWireDelay	(SBDATI1_ipd,SBDATI1,tipd_SBDATI1);
VitalWireDelay	(SBDATI0_ipd,SBDATI0,tipd_SBDATI0);
VitalWireDelay	(MI_ipd,MI,tipd_MI);
VitalWireDelay	(SI_ipd,SI,tipd_SI);
VitalWireDelay	(SCKI_ipd,SCKI,tipd_SCKI);
VitalWireDelay	(SCSNI_ipd,SCSNI,tipd_SCSNI);
End block;
----------------------------------------------------------------------
-- BEHAVIOR SECTION
----------------------------------------------------------------------

spiU:SB_SPI_CORE
generic map (
                  BUS_ADDR74 => BUS_ADDR74 
         )         
Port map(

	   SBDATO7   => SBDATO7_zd,  
      SBDATO6  => SBDATO6_zd, 
      SBDATO5   => SBDATO5_zd,  
      SBDATO4   => SBDATO4_zd,  
      SBDATO3   => SBDATO3_zd,  
      SBDATO2   => SBDATO2_zd,  
      SBDATO1   => SBDATO1_zd,  
      SBDATO0   => SBDATO0_zd,  
      SBACKO   => SBACKO_zd,  
      SPIIRQ   => SPIIRQ_zd,  
      SPIWKUP   => SPIWKUP_zd,  
      SO   => SO_zd,  
      SOE   => SOE_zd,  
      MO   => MO_zd,  
      MOE   => MOE_zd,  
	   SCKO => SCKO_zd,
		SCKOE => SCKOE_zd,
		MCSNO3 => MCSNO3_zd,
		MCSNO2 => MCSNO2_zd,
		MCSNO1 => MCSNO1_zd,
		MCSNO0 => MCSNO0_zd,
		MCSNOE3 => MCSNOE3_zd,
		MCSNOE2 => MCSNOE2_zd,
		MCSNOE1 => MCSNOE1_zd,
		MCSNOE0 => MCSNOE0_zd,
	
		SBCLKI => SBCLKI_ipd,
		SBRWI => SBRWI_ipd,
		SBSTBI => SBSTBI_ipd,
		SBADRI7 => SBADRI7_ipd,
		SBADRI6 => SBADRI6_ipd,
		SBADRI5 => SBADRI5_ipd,
		SBADRI4 => SBADRI4_ipd,
		SBADRI3 => SBADRI3_ipd,
		SBADRI2 => SBADRI2_ipd,
		SBADRI1 => SBADRI1_ipd,
		SBADRI0 => SBADRI0_ipd,
		SBDATI7 => SBDATI7_ipd,
		SBDATI6 => SBDATI6_ipd,
		SBDATI5 => SBDATI5_ipd,
		SBDATI4 => SBDATI4_ipd,
		SBDATI3 => SBDATI3_ipd,
		SBDATI2 => SBDATI2_ipd,
		SBDATI1 => SBDATI1_ipd,
		SBDATI0 => SBDATI0_ipd,
		MI => MI_ipd,
		SI => SI_ipd,
		SCKI => SCKI_ipd,
		SCSNI => SCSNI_ipd

);
	
-------------------------------------------------------------------
--VITAL timing check
------------------------------------------------------------------
VITALTimingCheck : process (SBCLKI_ipd, SBRWI_ipd, SBSTBI_ipd, SBADRI7_ipd, SBADRI6_ipd, SBADRI5_ipd, SBADRI4_ipd, SBADRI3_ipd, SBADRI2_ipd, SBADRI1_ipd, SBADRI0_ipd, SBDATI7_ipd, SBDATI6_ipd, SBDATI5_ipd, SBDATI4_ipd, SBDATI3_ipd, SBDATI2_ipd, SBDATI1_ipd, SBDATI0_ipd, MI_ipd, SI_ipd,SCKI_ipd,SCSNI_ipd)

    variable Tviol_SBRWI_SBCLKI_posedge      : std_ulogic := '0';
    variable Tviol_SBSTBI_SBCLKI_posedge     : std_ulogic := '0';
    variable Tviol_SCLI_SBCLKI_posedge       : std_ulogic := '0';
    variable Tviol_SDATI_SBCLKI_posedge      : std_ulogic := '0';
    variable Tviol_SBADRI7_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBADRI6_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBADRI5_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBADRI4_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBADRI3_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBADRI2_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBADRI1_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBADRI0_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBDATI7_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBDATI6_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBDATI5_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBDATI4_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBDATI3_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBDATI2_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBDATI1_SBCLKI_posedge    : std_ulogic := '0';
    variable Tviol_SBDATI0_SBCLKI_posedge    : std_ulogic := '0';
  	variable Tviol_MI_SCKO_posedge    		 : std_ulogic := '0';
	variable Tviol_SI_SCKI_posedge     		 : std_ulogic := '0';
	variable Tviol_SCSNI_SCKI_posedge     	 : std_ulogic := '0';	
	----------------------------added----------------------------
	variable Tviol_MI_SCKO_negedge    		 : std_ulogic := '0';
	variable Tviol_SI_SCKI_negedge     		 : std_ulogic := '0';
	variable Tviol_SCSNI_SCKI_negedge     	 : std_ulogic := '0';
	-------------------------------------------------------------

	variable Tmkr_SBRWI_SBCLKI_posedge       : VitalTimingDataType := VitalTimingDataInit;
    variable Tmkr_SBSTBI_SBCLKI_posedge      : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_SBRWI_SCLI_posedge     	 : VitalTimingDataType := VitalTimingDataInit;
    variable Tmkr_SDATI_SBCLKI_posedge       : VitalTimingDataType := VitalTimingDataInit;
    variable Tmkr_SBADRI7_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
    variable Tmkr_SBADRI6_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
    variable Tmkr_SBADRI5_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_SBADRI4_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
    variable Tmkr_SBADRI3_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
    variable Tmkr_SBADRI2_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
    variable Tmkr_SBADRI1_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
    variable Tmkr_SBADRI0_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_SBDATI7_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
    variable Tmkr_SBDATI6_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
    variable Tmkr_SBDATI5_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_SBDATI4_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
    variable Tmkr_SBDATI3_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
    variable Tmkr_SBDATI2_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
    variable Tmkr_SBDATI1_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
    variable Tmkr_SBDATI0_SBCLKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MI_SCKO_posedge     : VitalTimingDataType := VitalTimingDataInit;		  
	variable Tmkr_SI_SCKI_posedge     : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_SCSNI_SCKI_posedge     : VitalTimingDataType := VitalTimingDataInit; 
	----------------------------added---------------------------- 
	variable Tmkr_MI_SCKO_negedge    		 : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_SI_SCKI_negedge     		 : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_SCSNI_SCKI_negedge     	 : VitalTimingDataType := VitalTimingDataInit;
	-------------------------------------------------------------


begin
if (TimingChecksOn) then
      VitalSetupHoldCheck (
        Violation      => Tviol_SBRWI_SBCLKI_posedge,
        TimingData     => Tmkr_SBRWI_SBCLKI_posedge,
        TestSignal     => SBRWI_ipd,
        TestSignalName => "SBRWI",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBRWI_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBRWI_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBRWI_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBRWI_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_SPI",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);
 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBSTBI_SBCLKI_posedge,
        TimingData     => Tmkr_SBSTBI_SBCLKI_posedge,
        TestSignal     => SBSTBI_ipd,
        TestSignalName => "SBSTBI",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBSTBI_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBSTBI_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBSTBI_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBSTBI_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_SPI",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);
  		 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBADRI7_SBCLKI_posedge,
        TimingData     => Tmkr_SBADRI7_SBCLKI_posedge,
        TestSignal     => SBADRI7_ipd,
        TestSignalName => "SBADRI7",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBADRI7_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBADRI7_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBADRI7_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBADRI7_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_SPI",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);		
 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBADRI6_SBCLKI_posedge,
        TimingData     => Tmkr_SBADRI6_SBCLKI_posedge,
        TestSignal     => SBADRI6_ipd,
        TestSignalName => "SBADRI6",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBADRI6_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBADRI6_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBADRI6_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBADRI6_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_SPI",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);		

		 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBADRI5_SBCLKI_posedge,
        TimingData     => Tmkr_SBADRI5_SBCLKI_posedge,
        TestSignal     => SBADRI5_ipd,
        TestSignalName => "SBADRI5",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBADRI5_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBADRI5_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBADRI5_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBADRI5_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_SPI",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);		
		
 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBADRI4_SBCLKI_posedge,
        TimingData     => Tmkr_SBADRI4_SBCLKI_posedge,
        TestSignal     => SBADRI4_ipd,
        TestSignalName => "SBADRI4",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBADRI4_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBADRI4_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBADRI4_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBADRI4_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_SPI",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);	
 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBADRI3_SBCLKI_posedge,
        TimingData     => Tmkr_SBADRI3_SBCLKI_posedge,
        TestSignal     => SBADRI3_ipd,
        TestSignalName => "SBADRI3",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBADRI3_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBADRI3_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBADRI3_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBADRI3_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_SPI",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);		
 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBADRI2_SBCLKI_posedge,
        TimingData     => Tmkr_SBADRI2_SBCLKI_posedge,
        TestSignal     => SBADRI2_ipd,
        TestSignalName => "SBADRI2",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBADRI2_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBADRI2_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBADRI2_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBADRI2_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_SPI",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);
 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBADRI1_SBCLKI_posedge,
        TimingData     => Tmkr_SBADRI1_SBCLKI_posedge,
        TestSignal     => SBADRI1_ipd,
        TestSignalName => "SBADRI1",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBADRI1_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBADRI1_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBADRI1_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBADRI1_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_SPI",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);	
 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBADRI0_SBCLKI_posedge,
        TimingData     => Tmkr_SBADRI0_SBCLKI_posedge,
        TestSignal     => SBADRI0_ipd,
        TestSignalName => "SBADRI0",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBADRI0_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBADRI0_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBADRI0_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBADRI0_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_SPI",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);	
	

	
		 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBDATI7_SBCLKI_posedge,
        TimingData     => Tmkr_SBDATI7_SBCLKI_posedge,
        TestSignal     => SBDATI7_ipd,
        TestSignalName => "SBDATI7",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBDATI7_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBDATI7_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBDATI7_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBDATI7_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_SPI",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);		
 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBDATI6_SBCLKI_posedge,
        TimingData     => Tmkr_SBDATI6_SBCLKI_posedge,
        TestSignal     => SBDATI6_ipd,
        TestSignalName => "SBDATI6",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBDATI6_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBDATI6_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBDATI6_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBDATI6_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_SPI",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);		

		 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBDATI5_SBCLKI_posedge,
        TimingData     => Tmkr_SBDATI5_SBCLKI_posedge,
        TestSignal     => SBDATI5_ipd,
        TestSignalName => "SBDATI5",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBDATI5_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBDATI5_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBDATI5_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBDATI5_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_SPI",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);		
		
 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBDATI4_SBCLKI_posedge,
        TimingData     => Tmkr_SBDATI4_SBCLKI_posedge,
        TestSignal     => SBDATI4_ipd,
        TestSignalName => "SBDATI4",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBDATI4_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBDATI4_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBDATI4_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBDATI4_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_SPI",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);	
 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBDATI3_SBCLKI_posedge,
        TimingData     => Tmkr_SBDATI3_SBCLKI_posedge,
        TestSignal     => SBDATI3_ipd,
        TestSignalName => "SBDATI3",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBDATI3_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBDATI3_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBDATI3_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBDATI3_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_SPI",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);		
 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBDATI2_SBCLKI_posedge,
        TimingData     => Tmkr_SBDATI2_SBCLKI_posedge,
        TestSignal     => SBDATI2_ipd,
        TestSignalName => "SBDATI2",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBDATI2_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBDATI2_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBDATI2_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBDATI2_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_SPI",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);
 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBDATI1_SBCLKI_posedge,
        TimingData     => Tmkr_SBDATI1_SBCLKI_posedge,
        TestSignal     => SBDATI1_ipd,
        TestSignalName => "SBDATI1",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBDATI1_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBDATI1_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBDATI1_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBDATI1_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_SPI",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);	
 
      VitalSetupHoldCheck (
        Violation      => Tviol_SBDATI0_SBCLKI_posedge,
        TimingData     => Tmkr_SBDATI0_SBCLKI_posedge,
        TestSignal     => SBDATI0_ipd,
        TestSignalName => "SBDATI0",
        RefSignal      => SBCLKI_ipd,
        RefSignalName  => "SBCLKI",
        SetupHigh      => tsetup_SBDATI0_SBCLKI_posedge_posedge,
        SetupLow       => tsetup_SBDATI0_SBCLKI_negedge_posedge,
        HoldLow        => thold_SBDATI0_SBCLKI_negedge_posedge,
        HoldHigh       => thold_SBDATI0_SBCLKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_SPI",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);	
		
	
		VitalSetupHoldCheck (
        Violation      => Tviol_MI_SCKO_posedge,
        TimingData     => Tmkr_MI_SCKO_posedge,
        TestSignal     => MI,
        TestSignalName => "MI",
      	RefSignal      => SCKO_zd,
        RefSignalName  => "SCKO",
        SetupHigh      => tsetup_MI_SCKO_posedge_posedge,
        SetupLow       => tsetup_MI_SCKO_negedge_posedge,
        HoldLow        => thold_MI_SCKO_negedge_posedge,
        HoldHigh       => thold_MI_SCKO_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_SPI",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);
	VitalSetupHoldCheck (
        Violation      => Tviol_SI_SCKI_posedge,
        TimingData     => Tmkr_SI_SCKI_posedge,
        TestSignal     => SI_ipd,
        TestSignalName => "SI",
        RefSignal      => SCKI_ipd,
        RefSignalName  => "SCKI",
        SetupHigh      => tsetup_SI_SCKI_posedge_posedge,
        SetupLow       => tsetup_SI_SCKI_negedge_posedge,
        HoldLow        => thold_SI_SCKI_negedge_posedge,
        HoldHigh       => thold_SI_SCKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_SPI",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);	
	VitalSetupHoldCheck (
        Violation      => Tviol_SCSNI_SCKI_posedge,
        TimingData     => Tmkr_SCSNI_SCKI_posedge,
        TestSignal     => SCSNI_ipd,
        TestsignalName => "SCSNI",
        RefSignal      => SCKI_ipd,
        RefSignalName  => "SCKI",
        SetupHigh      => tsetup_SCSNI_SCKI_posedge_posedge,
        SetupLow       => tsetup_SCSNI_SCKI_negedge_posedge,
        HoldLow        => thold_SCSNI_SCKI_negedge_posedge,
        HoldHigh       => thold_SCSNI_SCKI_posedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_SPI",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);	
		
		------------------------added--------------------
	VitalSetupHoldCheck (
        Violation      => Tviol_MI_SCKO_negedge,
        TimingData     => Tmkr_MI_SCKO_negedge,
        TestSignal     => MI,
        TestSignalName => "MI",
      	RefSignal      => SCKO_zd,
        RefSignalName  => "SCKO",
        SetupHigh      => tsetup_MI_SCKO_posedge_negedge,
        SetupLow       => tsetup_MI_SCKO_negedge_negedge,
        HoldLow        => thold_MI_SCKO_negedge_negedge,
        HoldHigh       => thold_MI_SCKO_posedge_negedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_SPI",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);
	VitalSetupHoldCheck (
        Violation      => Tviol_SI_SCKI_negedge,
        TimingData     => Tmkr_SI_SCKI_negedge,
        TestSignal     => SI_ipd,
        TestSignalName => "SI",
        RefSignal      => SCKI_ipd,
        RefSignalName  => "SCKI",
        SetupHigh      => tsetup_SI_SCKI_posedge_negedge,
        SetupLow       => tsetup_SI_SCKI_negedge_negedge,
        HoldLow        => thold_SI_SCKI_negedge_negedge,
        HoldHigh       => thold_SI_SCKI_posedge_negedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_SPI",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);	
	VitalSetupHoldCheck (
        Violation      => Tviol_SCSNI_SCKI_negedge,
        TimingData     => Tmkr_SCSNI_SCKI_negedge,
        TestSignal     => SCSNI_ipd,
        TestsignalName => "SCSNI",
        RefSignal      => SCKI_ipd,
        RefSignalName  => "SCKI",
        SetupHigh      => tsetup_SCSNI_SCKI_posedge_negedge,
        SetupLow       => tsetup_SCSNI_SCKI_negedge_negedge,
        HoldLow        => thold_SCSNI_SCKI_negedge_negedge,
        HoldHigh       => thold_SCSNI_SCKI_posedge_negedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_SPI",
        Xon            => Xon,
        MsgOn          => true,
        MsgSeverity    => warning);	
		-------------------------------------------------

end if;
end process VITALTimingCheck;




 




VITALPathDelay0: process (SBCLKI_ipd,SBDATO0_zd,SBDATO1_zd,SBDATO2_zd,SBDATO3_zd,SBDATO4_zd,SBDATO5_zd,SBDATO6_zd,SBDATO7_zd)
		
variable SBDATO7_GlitchData : VitalGlitchDataType; 
variable SBDATO6_GlitchData : VitalGlitchDataType; 
variable SBDATO5_GlitchData : VitalGlitchDataType;
variable SBDATO4_GlitchData : VitalGlitchDataType;
variable SBDATO3_GlitchData : VitalGlitchDataType;
variable SBDATO2_GlitchData : VitalGlitchDataType;
variable SBDATO1_GlitchData : VitalGlitchDataType;
variable SBDATO0_GlitchData : VitalGlitchDataType;

variable        SBDATO7_tmp  : std_ulogic := 'X';
variable        SBDATO6_tmp  : std_ulogic := 'X';
variable        SBDATO5_tmp  : std_ulogic := 'X';
variable        SBDATO4_tmp  : std_ulogic := 'X';
variable        SBDATO3_tmp  : std_ulogic := 'X';
variable        SBDATO2_tmp  : std_ulogic := 'X';
variable        SBDATO1_tmp  : std_ulogic := 'X';
variable        SBDATO0_tmp  : std_ulogic := 'X';

begin	 
	SBDATO7_tmp:=SBDATO7_zd;	
	SBDATO6_tmp:=SBDATO6_zd;
	SBDATO5_tmp:=SBDATO5_zd;
	SBDATO4_tmp:=SBDATO4_zd;
	SBDATO3_tmp:=SBDATO3_zd;
	SBDATO2_tmp:=SBDATO2_zd;
	SBDATO1_tmp:=SBDATO1_zd;  
	SBDATO0_tmp:=SBDATO0_zd;
  VitalPathDelay01 (
      OutSignal                 => SBDATO7,
      GlitchData                => SBDATO7_GlitchData,
      OutSignalName             => "SBDATO7",
      OutTemp                   => SBDATO7_tmp,
      Paths                     => (0 => (SBCLKI_ipd'last_event, tpd_SBCLKI_SBDATO7_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);	
	  
	
VitalPathDelay01 (
      OutSignal                 => SBDATO6,
      GlitchData                => SBDATO6_GlitchData,
      OutSignalName             => "SBDATO6",
      OutTemp                   => SBDATO6_tmp,
      Paths                     => (0 => (SBCLKI_ipd'last_event, tpd_SBCLKI_SBDATO6_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

	
  VitalPathDelay01 (
      OutSignal                 => SBDATO5,
      GlitchData                => SBDATO5_GlitchData,
      OutSignalName             => "SBDATO5",
      OutTemp                   => SBDATO5_tmp,
      Paths                     => (0 => (SBCLKI_ipd'last_event, tpd_SBCLKI_SBDATO5_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

  VitalPathDelay01 (
      OutSignal                 => SBDATO4,
      GlitchData                => SBDATO4_GlitchData,
      OutSignalName             => "SBDATO4",
      OutTemp                   => SBDATO4_tmp,
      Paths                     => (0 => (SBCLKI_ipd'last_event, tpd_SBCLKI_SBDATO4_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
	
  VitalPathDelay01 (
      OutSignal                 => SBDATO3,
      GlitchData                => SBDATO3_GlitchData,
      OutSignalName             => "SBDATO3",
      OutTemp                   => SBDATO3_tmp,
      Paths                     => (0 => (InputChangeTime=>SBCLKI_ipd'last_event,
	  PathDelay=>tpd_SBCLKI_SBDATO3_posedge,
	  PathCondition=>true)	),
     Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning
	  );

	
  VitalPathDelay01 (
      OutSignal                 => SBDATO2,
      GlitchData                => SBDATO2_GlitchData,
      OutSignalName             => "SBDATO2",
      OutTemp                   => SBDATO2_tmp,
      Paths                     => (0 => (SBCLKI_ipd'last_event, tpd_SBCLKI_SBDATO2_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
	
	
  VitalPathDelay01 (
      OutSignal                 => SBDATO1,
      GlitchData                => SBDATO1_GlitchData,
      OutSignalName             => "SBDATO1",
      OutTemp                   => SBDATO1_tmp,
      Paths                     => (0 => (SBCLKI_ipd'last_event, tpd_SBCLKI_SBDATO1_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
	
  VitalPathDelay01 (
      OutSignal                 => SBDATO0,
      GlitchData                => SBDATO0_GlitchData,
      OutSignalName             => "SBDATO0",
      OutTemp                   => SBDATO0_tmp,
      Paths                     => (0 => (SBCLKI_ipd'last_event, tpd_SBCLKI_SBDATO0_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
 
	end process VITALPathDelay0;  
	
	
VITALPathDelay   : process (SBCLKI_ipd,SBACKO_zd,SCKO_zd,SPIIRQ_zd, SOE_zd,SO_zd, MCSNOE0_zd,MCSNOE1_zd,MCSNOE2_zd,MCSNOE3_zd,MCSNO0_zd,MCSNO1_zd,MCSNO2_zd,MCSNO3_zd,MOE_zd,MO_zd,SPIWKUP_zd)
variable SBACKO_GlitchData : VitalGlitchDataType;
variable SPIIRQ_GlitchData : VitalGlitchDataType;
variable SPIWKUP_GlitchData : VitalGlitchDataType;
variable SO_GlitchData : VitalGlitchDataType;
variable SOE_GlitchData : VitalGlitchDataType;
variable MO_GlitchData : VitalGlitchDataType;
variable MOE_GlitchData : VitalGlitchDataType;
variable SCKO_GlitchData : VitalGlitchDataType;
variable SCKOE_GlitchData : VitalGlitchDataType;
variable MCSNO3_GlitchData : VitalGlitchDataType;
variable MCSNO2_GlitchData : VitalGlitchDataType;
variable MCSNO1_GlitchData : VitalGlitchDataType;
variable MCSNO0_GlitchData : VitalGlitchDataType;
variable MCSNOE3_GlitchData : VitalGlitchDataType;
variable MCSNOE2_GlitchData : VitalGlitchDataType;
variable MCSNOE1_GlitchData : VitalGlitchDataType;
variable MCSNOE0_GlitchData : VitalGlitchDataType;	  


variable        SBACKO_tmp  : std_ulogic := 'X';
variable        SPIIRQ_tmp  : std_ulogic := 'X';
variable        SPIWKUP_tmp  : std_ulogic := 'X';
variable        SO_tmp  : std_ulogic := 'X';
variable        SOE_tmp  : std_ulogic := 'X';
variable        MO_tmp  : std_ulogic := 'X';
variable        MOE_tmp  : std_ulogic := 'X';
variable        SCKO_tmp  : std_ulogic := 'X';
variable        SCKOE_tmp  : std_ulogic := 'X';
variable        MCSNO3_tmp  : std_ulogic := 'X';
variable        MCSNO2_tmp  : std_ulogic := 'X';
variable        MCSNO1_tmp  : std_ulogic := 'X';
variable        MCSNO0_tmp  : std_ulogic := 'X';
variable        MCSNOE3_tmp  : std_ulogic := 'X';
variable        MCSNOE2_tmp  : std_ulogic := 'X';
variable        MCSNOE1_tmp  : std_ulogic := 'X';
variable        MCSNOE0_tmp  : std_ulogic := 'X';

begin		   
	        SBACKO_tmp := SBACKO_zd;
        SPIIRQ_tmp := SPIIRQ_zd;
        SPIWKUP_tmp := SPIWKUP_zd;
        SO_tmp := SO_zd;
        SOE_tmp := SOE_zd;
        MO_tmp := MO_zd;
        MOE_tmp := MOE_zd;
        SCKO_tmp := SCKO_zd;
        SCKOE_tmp := SCKOE_zd;
        MCSNO3_tmp := MCSNO3_zd;
        MCSNO2_tmp := MCSNO2_zd;
        MCSNO1_tmp := MCSNO1_zd;
        MCSNO0_tmp := MCSNO0_zd;
        MCSNOE3_tmp := MCSNOE3_zd;
        MCSNOE2_tmp := MCSNOE2_zd;
        MCSNOE1_tmp := MCSNOE1_zd;
        MCSNOE0_tmp := MCSNOE0_zd;
  VitalPathDelay01 (
      OutSignal                 => SBACKO,
      GlitchData                => SBACKO_GlitchData,
      OutSignalName             => "SBACKO",
      OutTemp                   => SBACKO_tmp,
      Paths                     => (0 => (SBCLKI_ipd'last_event, tpd_SBCLKI_SBACKO_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning); 
	


	 
VitalPathDelay01 (
      OutSignal                 => SPIIRQ,
      GlitchData                => SPIIRQ_GlitchData,
      OutSignalName             => "SPIIRQ",
      OutTemp                   => SPIIRQ_tmp,
      Paths                     => (0 => (SBCLKI_ipd'last_event, tpd_SBCLKI_SPIIRQ_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);		   

	  
	  VitalPathDelay01 (
      OutSignal                 => SPIWKUP,
      GlitchData                => SPIWKUP_GlitchData,
      OutSignalName             => "SPIWKUP",
      OutTemp                   => SPIWKUP_tmp,
      Paths                     => (0 => (SBCLKI_ipd'last_event, tpd_SBCLKI_SPIWKUP_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);		   
	  


VitalPathDelay01 (
      OutSignal                 => MO,
      GlitchData                => MO_GlitchData,
      OutSignalName             => "MO",
      OutTemp                   => MO_tmp,
      Paths                     => (0 => (SCKO_zd'last_event, tpd_SCKO_MO_posedge, true)	),	 
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

	  
  
VitalPathDelay01 (
      OutSignal                 => MO,
      GlitchData                => MO_GlitchData,
      OutSignalName             => "MO",
      OutTemp                   => MO_tmp,
      Paths                     => (0 => (SCKO_zd'last_event, tpd_SCKO_MO_negedge, true)	),	 
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
	  


VitalPathDelay01 (
      OutSignal                 => MOE,
      GlitchData                => MOE_GlitchData,
      OutSignalName             => "MOE",
      OutTemp                   => MOE_tmp,
      Paths                     => (0 => (SCKO_zd'last_event, tpd_SCKO_MOE_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
	  
	  

VitalPathDelay01 (
      OutSignal                 => MCSNO3,
      GlitchData                => MCSNO3_GlitchData,
      OutSignalName             => "MCSNO3",
      OutTemp                   => MCSNO3_tmp,
      Paths                     => (0 => (SCKO_zd'last_event, tpd_SCKO_MCSNO3_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

	  

VitalPathDelay01 (
      OutSignal                 => MCSNO2,
      GlitchData                => MCSNO2_GlitchData,
      OutSignalName             => "MCSNO2",
      OutTemp                   => MCSNO2_tmp,
      Paths                     => (0 => (SCKO_zd'last_event, tpd_SCKO_MCSNO2_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
	  

VitalPathDelay01 (
      OutSignal                 => MCSNO1,
      GlitchData                => MCSNO1_GlitchData,
      OutSignalName             => "MCSNO1",
      OutTemp                   => MCSNO1_tmp,
      Paths                     => (0 => (SCKO_zd'last_event, tpd_SCKO_MCSNO1_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
	  

VitalPathDelay01 (
      OutSignal                 => MCSNO0,
      GlitchData                => MCSNO0_GlitchData,
      OutSignalName             => "MCSNO0",
      OutTemp                   => MCSNO0_tmp,
      Paths                     => (0 => (SCKO_zd'last_event, tpd_SCKO_MCSNO0_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
	  
	  

VitalPathDelay01 (
      OutSignal                 => MCSNOE3,
      GlitchData                => MCSNOE3_GlitchData,
      OutSignalName             => "MCSNOE3",
      OutTemp                   => MCSNOE3_tmp,
      Paths                     => (0 => (SCKO_zd'last_event, tpd_SCKO_MCSNOE3_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
	  
	  

VitalPathDelay01 (
      OutSignal                 => MCSNOE2,
      GlitchData                => MCSNOE2_GlitchData,
      OutSignalName             => "MCSNOE2",
      OutTemp                   => MCSNOE2_tmp,
      Paths                     => (0 => (SCKO_zd'last_event, tpd_SCKO_MCSNOE2_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
	  
	  

VitalPathDelay01 (
      OutSignal                 => MCSNOE1,
      GlitchData                => MCSNOE1_GlitchData,
      OutSignalName             => "MCSNOE1",
      OutTemp                   => MCSNOE1_tmp,
      Paths                     => (0 => (SCKO_zd'last_event, tpd_SCKO_MCSNOE1_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
	  
	  

VitalPathDelay01 (
      OutSignal                 => MCSNOE0,
      GlitchData                => MCSNOE0_GlitchData,
      OutSignalName             => "MCSNOE0",
      OutTemp                   => MCSNOE0_tmp,
      Paths                     => (0 => (SCKO_zd'last_event, tpd_SCKO_MCSNOE0_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);		   
	  

VitalPathDelay01 (
      OutSignal                 => SO,
      GlitchData                => SO_GlitchData,
      OutSignalName             => "SO",
      OutTemp                   => SO_tmp,
      Paths                     => (0 => (SCKI_ipd'last_event, tpd_SCKI_SO_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);	 
	  
	  

VitalPathDelay01 (
      OutSignal                 => SO,
      GlitchData                => SO_GlitchData,
      OutSignalName             => "SO",
      OutTemp                   => SO_tmp,
      Paths                     => (0 => (SCKI_ipd'last_event, tpd_SCKI_SO_negedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
	  
	  

VitalPathDelay01 (	   	

      OutSignal                 => SOE,
      GlitchData                => SOE_GlitchData,
      OutSignalName             => "SOE",
      OutTemp                   => SOE_tmp,
      Paths                     => (0 => (SCKI_ipd'last_event, tpd_SCKI_SOE_posedge, true)	),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);  

  end process VITALPathDelay;

end SB_SPI_V;


-------------------------------------------------
---     	SB_LSOSC 		-------
------------------------------------------------
library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use IEEE.Vital_Primitives.all;
use IEEE.VITAL_Timing.all;
entity  SB_LSOSC  is 
	generic(
	Xon   : boolean := true;
    	MsgOn : boolean := true;

	tipd_ENACLKK: VitalDelayType01 := (0.000 ns, 0.000 ns);
      	tpd_ENACLKK_CLKK : VitalDelayType01 := (0.000 ns, 0.000 ns)
 ); 
port(
    CLKK : out std_logic;
    ENACLKK : in std_logic
    );
 attribute VITAL_LEVEL0 of			    
    SB_LSOSC  : entity is true;
end SB_LSOSC ;

architecture SB_LSOSC_V of SB_LSOSC is
  attribute VITAL_LEVEL0 of
    SB_LSOSC_V : architecture is true;

signal ENACLKK_ipd: std_ulogic := 'X';
signal CLKK_zd  : std_ulogic	:='X'; 

component SB_LSOSC_CORE
port (
	ENACLKK : IN std_logic;
	CLKK : OUT std_logic
);
end component;
			  

begin
  WireDelay : block
  begin
    VitalWireDelay (ENACLKK_ipd, ENACLKK, tipd_ENACLKK);
  end block;
----------------------------------------------------------------
-- BEHAVIOR SECTION
----------------------------------------------------------------
LS: SB_LSOSC_CORE
port map(
	ENACLKK=> ENACLKK_ipd,
	CLKK=> CLKK_zd
		);
VITALPathDelay :process (ENACLKK_ipd,CLKK_zd)
variable CLKK_GlitchData : VitalGlitchDataType;		  
variable CLKK_tmp:std_ulogic:='X';
begin			 
	CLKK_tmp:=CLKK_zd;
VitalPathDelay01 (
      OutSignal                 => CLKK,
      GlitchData                => CLKK_GlitchData,
      OutSignalName             => "CLKK",
      OutTemp                   => CLKK_tmp,
      Paths                     => (0 =>(ENACLKK_ipd'last_event, tpd_ENACLKK_CLKK, true)),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
end process;
end 	SB_LSOSC_V; 

--------------------------------------------------------------
---     	SB_HSOSC 		-------
------------------------------------------------

library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use IEEE.Vital_Primitives.all;
use IEEE.VITAL_Timing.all;
entity  SB_HSOSC  is 
	generic(
	Xon   : boolean := true;
    MsgOn : boolean := true;

	tipd_ENACLKM: VitalDelayType01 := (0.000 ns, 0.000 ns);
    tpd_ENACLKM_CLKM : VitalDelayType01 := (0.000 ns, 0.000 ns)
 ); 
port(
    CLKM : out std_logic;
    ENACLKM : in std_logic
    );
 attribute VITAL_LEVEL0 of
    SB_HSOSC  : entity is true;			    
end SB_HSOSC ;

architecture SB_HSOSC_V of SB_HSOSC is
  attribute VITAL_LEVEL0 of
    SB_HSOSC_V : architecture is true;

signal ENACLKM_ipd: std_ulogic 	:= 'X';
signal CLKM_zd   :   std_ulogic	:='X';

component SB_HSOSC_CORE
port (
	ENACLKM : IN std_logic;
	CLKM : OUT std_logic
);
end component;

begin
--wire delay
  WireDelay : block
  begin
    VitalWireDelay (ENACLKM_ipd, ENACLKM, tipd_ENACLKM);
  end block;

----------------------------------------------------------------
-- BEHAVIOR SECTION
----------------------------------------------------------------
HS: SB_HSOSC_CORE
port map(
	ENACLKM=> ENACLKM_ipd,
	CLKM=> CLKM_zd
		);

-- PATH DELAY
VITALPathDelay :process (ENACLKM_ipd,CLKM_zd)
variable CLKM_GlitchData : VitalGlitchDataType;	 
variable CLKM_tmp :std_ulogic:='X';
begin							   
	CLKM_tmp:=CLKM_zd;
VitalPathDelay01 (
      OutSignal                 => CLKM,
      GlitchData                => CLKM_GlitchData,
      OutSignalName             => "CLKM",
      OutTemp                   => CLKM_tmp,
      Paths                     => (0 =>(ENACLKM_ipd'last_event, tpd_ENACLKM_CLKM, true)),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
end process;
end 	SB_HSOSC_V; 

-- ICE5LP Primitives 

------------------------------------------------
---     	SB_IO_OD 		-------
------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
--library	work;
use IEEE.Vital_Primitives.all;
use IEEE.VITAL_Timing.all;
use	work.std_logic_SBT.all;

entity	SB_IO_OD is

	generic (
			TimingChecksOn : boolean := true;
			Xon   : boolean := true;
			MsgOn : boolean := true;
			tipd_DOUT1: VitalDelayType01 := (0.000 ns, 0.000 ns);
			tipd_DOUT0: VitalDelayType01 := (0.000 ns, 0.000 ns);
			tipd_CLOCKENABLE: VitalDelayType01 := (0.000 ns, 0.000 ns);
			tipd_LATCHINPUTVALUE: VitalDelayType01 := (0.000 ns, 0.000 ns);
			tipd_INPUTCLK: VitalDelayType01 := (0.000 ns, 0.000 ns);
			tipd_OUTPUTENABLE: VitalDelayType01 := (0.000 ns, 0.000 ns);
			tipd_OUTPUTCLK: VitalDelayType01 := (0.000 ns, 0.000 ns);
			tipd_PACKAGEPIN: VitalDelayType01 := (0.000 ns, 0.000 ns);
			
			tpd_PACKAGEPIN_DIN0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
			tpd_PACKAGEPIN_DIN1  : VitalDelayType01 := (0.000 ns, 0.000 ns);
			tpd_INPUTCLK_DIN0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
			tpd_INPUTCLK_DIN1  : VitalDelayType01 := (0.000 ns, 0.000 ns);
			tpd_DOUT0_PACKAGEPIN : VitalDelayType01 := (0.000 ns, 0.000 ns);
			tpd_DOUT1_PACKAGEPIN : VitalDelayType01 := (0.000 ns, 0.000 ns);
			tpd_OUTPUTENABLE_PACKAGEPIN : VitalDelayType01 := (0.000 ns, 0.000 ns);
			tpd_INPUTCLK_PACKAGEPIN : VitalDelayType01 := (0.000 ns, 0.000 ns);
			tpd_OUTPUTCLK_PACKAGEPIN  : VitalDelayType01 := (0.000 ns, 0.000 ns);
			tpd_LATCHINPUTVALUE_DIN1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
			tpd_LATCHINPUTVALUE_DIN0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
			tpd_INPUTCLK_DIN0_posedge 			: VitalDelayType01 := (0.000 ns, 0.000 ns);
            tpd_INPUTCLK_DIN1_negedge 			: VitalDelayType01 := (0.000 ns, 0.000 ns);	
			tpd_OUTPUTCLK_PACKAGEPIN_posedge 		: VitalDelayType01 := (0.000 ns, 0.000 ns);
			tpd_OUTPUTCLK_PACKAGEPIN_negedge 		: VitalDelayType01 := (0.000 ns, 0.000 ns);
			
			tsetup_CLOCKENABLE_INPUTCLK_posedge_posedge  : VitalDelayType     := 0 ns;
			tsetup_CLOCKENABLE_INPUTCLK_negedge_posedge  : VitalDelayType     := 0 ns;
			tsetup_CLOCKENABLE_OUTPUTCLK_posedge_posedge  : VitalDelayType     := 0 ns;
			tsetup_CLOCKENABLE_OUTPUTCLK_negedge_posedge  : VitalDelayType     := 0 ns;
			tsetup_PACKAGEPIN_INPUTCLK_posedge_posedge  : VitalDelayType     := 0 ns;
			tsetup_PACKAGEPIN_INPUTCLK_negedge_posedge  : VitalDelayType     := 0 ns;
			tsetup_PACKAGEPIN_INPUTCLK_posedge_negedge  : VitalDelayType     := 0 ns;
			tsetup_PACKAGEPIN_INPUTCLK_negedge_negedge  : VitalDelayType     := 0 ns;
			tsetup_PACKAGEPIN_OUTPUTCLK_posedge_posedge  : VitalDelayType     := 0 ns;
			tsetup_PACKAGEPIN_OUTPUTCLK_negedge_posedge  : VitalDelayType     := 0 ns;
			tsetup_DOUT0_OUTPUTCLK_posedge_posedge  : VitalDelayType     := 0 ns;
			tsetup_DOUT0_OUTPUTCLK_negedge_posedge  : VitalDelayType     := 0 ns;
			tsetup_DOUT0_OUTPUTCLK_posedge_negedge  : VitalDelayType     := 0 ns;
			tsetup_DOUT0_OUTPUTCLK_negedge_negedgee  : VitalDelayType     := 0 ns;
			tsetup_DOUT1_OUTPUTCLK_posedge_posedge  : VitalDelayType     := 0 ns;
			tsetup_DOUT1_OUTPUTCLK_negedge_posedge  : VitalDelayType     := 0 ns;
			tsetup_DOUT1_OUTPUTCLK_posedge_negedge  : VitalDelayType     := 0 ns;
			tsetup_DOUT1_OUTPUTCLK_negedge_negedge  : VitalDelayType     := 0 ns;
			tsetup_OUTPUTENABLE_OUTPUTCLK_posedge_posedge  : VitalDelayType     := 0 ns;
			tsetup_OUTPUTENABLE_OUTPUTCLK_negedge_posedge  : VitalDelayType     := 0 ns;
			thold_CLOCKENABLE_INPUTCLK_posedge_posedge  : VitalDelayType     := 0 ns;
			thold_CLOCKENABLE_INPUTCLK_negedge_posedge  : VitalDelayType     := 0 ns;
			thold_CLOCKENABLE_OUTPUTCLK_posedge_posedge  : VitalDelayType     := 0 ns;
			thold_CLOCKENABLE_OUTPUTCLK_negedge_posedge  : VitalDelayType     := 0 ns;
			thold_PACKAGEPIN_INPUTCLK_posedge_posedge  : VitalDelayType     := 0 ns;
			thold_PACKAGEPIN_INPUTCLK_negedge_posedge  : VitalDelayType     := 0 ns;
			thold_PACKAGEPIN_INPUTCLK_posedge_negedge  : VitalDelayType     := 0 ns;
			thold_PACKAGEPIN_INPUTCLK_negedge_negedge  : VitalDelayType     := 0 ns;
			thold_PACKAGEPIN_OUTPUTCLK_posedge_posedge  : VitalDelayType     := 0 ns;
			thold_PACKAGEPIN_OUTPUTCLK_negedge_posedge  : VitalDelayType     := 0 ns;
			thold_DOUT0_OUTPUTCLK_posedge_posedge  : VitalDelayType     := 0 ns;
			thold_DOUT0_OUTPUTCLK_negedge_posedge  : VitalDelayType     := 0 ns;
			thold_DOUT0_OUTPUTCLK_posedge_negedge  : VitalDelayType     := 0 ns;
			thold_DOUT0_OUTPUTCLK_negedge_negedge  : VitalDelayType     := 0 ns;
			thold_DOUT1_OUTPUTCLK_posedge_posedge  : VitalDelayType     := 0 ns;
			thold_DOUT1_OUTPUTCLK_negedge_posedge  : VitalDelayType     := 0 ns;
			thold_DOUT1_OUTPUTCLK_posedge_negedge  : VitalDelayType     := 0 ns;
			thold_DOUT1_OUTPUTCLK_negedge_negedge  : VitalDelayType     := 0 ns;
			thold_OUTPUTENABLE_OUTPUTCLK_posedge_posedge  : VitalDelayType     := 0 ns;
			thold_OUTPUTENABLE_OUTPUTCLK_negedge_posedge  : VitalDelayType     := 0 ns;
			
			--tpd_ENACLKM_CLKM : VitalDelayType01 := (0.000 ns, 0.000 ns);
			NEG_TRIGGER : bit						:=	'0';
			PIN_TYPE	: bit_vector (5 downto 0)	:=	"000000"

			);
	port 
		(
		DOUT1 		    : in std_logic := 'L';
		DOUT0 		    : in std_logic := 'L';
		CLOCKENABLE		: in std_logic :='H';
		LATCHINPUTVALUE	: in std_logic;
		INPUTCLK			: in std_logic;
		
		DIN1				: out std_logic;
		DIN0				: out std_logic;
		OUTPUTENABLE		: in std_logic	:='H';
		OUTPUTCLK			: in std_logic;
		PACKAGEPIN			: inout	std_ulogic
		); 
				attribute VITAL_LEVEL0 of			    
    SB_IO_OD  : entity is true;
end SB_IO_OD ;

architecture SB_IO_OD_V of SB_IO_OD is
attribute VITAL_LEVEL0 of
    SB_IO_OD_V : architecture is true;
	signal DOUT1_ipd: std_ulogic := 'X';
	signal DOUT0_ipd: std_ulogic := 'X';
	signal CLOCKENABLE_ipd: std_ulogic := 'X';
	signal LATCHINPUTVALUE_ipd: std_ulogic := 'X';
	signal INPUTCLK_ipd: std_ulogic := 'X';
	signal OUTPUTENABLE_ipd: std_ulogic := 'X';
	signal OUTPUTCLK_ipd: std_ulogic := 'X';
	signal PACKAGEPIN_ipd: std_ulogic := 'X';
	
	signal DIN1_zd  : std_ulogic	:='X';
	signal DIN0_zd  : std_ulogic	:='X';
	signal PACKAGEPIN_zd  : std_ulogic	:='X';
	
	
	
	component	preio_physical
	port	(
			hold	:	in 	std_logic;
			rstio	:	in	std_logic;
			bs_en	:	in	std_logic;
			shift	:	in	std_logic;
			tclk	:	in	std_logic;
			inclk	:	in	std_logic;
			outclk	:	in	std_logic;
			update	:	in	std_logic;
			oepin	:	in	std_logic;
			sdi		:	in	std_logic;
			mode	:	in	std_logic;
			hiz_b	:	in	std_logic;
			sdo		:	out	std_logic;
			dout1	:	out	std_logic;
			dout0	:	out	std_logic;
			ddr1	:	in	std_logic;
			ddr0	:	in	std_logic;
			padin	:	in	std_logic;
			padout	:	out	std_logic;
			padoen	:	out	std_logic;
			cbit	:	in	std_logic_vector	(5 downto 0)
			);
	end component;

	signal	inclk_n, outclk_n, inclk, outclk,sdo	:	std_logic;
	
	signal	bs_en	:	std_logic	:='0';	--Boundary scan enable           
	signal	shift	:	std_logic	:='0';	--Boundary scan shift            
	signal	tclk	:	std_logic	:='0';	--Boundary scan clock            
	signal	update	:	std_logic	:='0';	--Boundary scan update           
	signal	sdi		:	std_logic	:='0';	--Boundary scan serial data in   
	signal	mode	:	std_logic	:='0';	--Boundary scan mode             
	signal	hiz_b	:	std_logic	:='1';	--Boundary scan Tristate control 
	
	signal	pin_cbit:	std_logic_vector(5 downto 0);
	signal	neg_trig:	std_logic;
	--signal	pull_up	:	std_logic;
	signal	hold,oepin,padoen,padout,padin	:	std_logic;
	signal INCLKE_sync , OUTCLKE_sync  	: std_logic;
begin

	WireDelay : block
  begin
    VitalWireDelay (DOUT1_ipd, DOUT1, tipd_DOUT1);
	VitalWireDelay (DOUT0_ipd, DOUT0, tipd_DOUT0);
	VitalWireDelay (CLOCKENABLE_ipd, CLOCKENABLE, tipd_CLOCKENABLE);
	VitalWireDelay (LATCHINPUTVALUE_ipd, LATCHINPUTVALUE, tipd_LATCHINPUTVALUE);
	VitalWireDelay (INPUTCLK_ipd, INPUTCLK, tipd_INPUTCLK);
	VitalWireDelay (OUTPUTENABLE_ipd, OUTPUTENABLE, tipd_OUTPUTENABLE);
	VitalWireDelay (OUTPUTCLK_ipd, OUTPUTCLK, tipd_OUTPUTCLK);
	VitalWireDelay (PACKAGEPIN_ipd, PACKAGEPIN, tipd_PACKAGEPIN);
	
  end block;
	
	pin_cbit	<=	TO_STDLOGICVECTOR	(PIN_TYPE);
	neg_trig	<=	TO_STDLOGIC	(NEG_TRIGGER);
	--pull_up		<=	TO_STDLOGIC	(PULLUP);

	inclk_n	<= 	INPUTCLK_ipd xor neg_trig;
	outclk_n<=	OUTPUTCLK_ipd xor neg_trig;
--	inclk	<=	inclk_n and CLOCK_ENABLE;
--	outclk	<=	outclk_n and CLOCK_ENABLE;

	process(inclk_n , CLOCKENABLE_ipd) is
         begin
                if(inclk_n ='0') then
                        INCLKE_sync  <= CLOCKENABLE_ipd;
                else
                        INCLKE_sync <= INCLKE_sync;
                end if ;
        end process;

        process(outclk_n , CLOCKENABLE_ipd) is
        begin
                if(outclk_n ='0') then
                        OUTCLKE_sync  <= CLOCKENABLE_ipd;
                else
                        OUTCLKE_sync <= OUTCLKE_sync;
                end if ;
        end process;

        inclk <= (inclk_n and INCLKE_sync);
        outclk <= (outclk_n and OUTCLKE_sync);
	
	hold	<=	LATCHINPUTVALUE_ipd;
	oepin	<=	OUTPUTENABLE_ipd;
	
	PACKAGE_PIN_i	:	process	(padoen, padout, PACKAGEPIN_ipd)
	begin
		padin	<=	PACKAGEPIN_ipd;
		if	((padoen='0')and (padout='0')) then
			PACKAGEPIN_zd	<=	'0';
		else
			PACKAGEPIN_zd	<=	'Z';
		end if;
	end process; 
-----------------------------------------------------------------	
	preio_physical_i	:	preio_physical
	port map	(
				hold	=>	hold,
				rstio	=>	'0',
				bs_en	=>	bs_en,
				shift	=>	shift,
				tclk	=>	tclk,
				inclk	=>	inclk,
				outclk	=>	outclk,
				update	=>	update,
				oepin	=>	oepin,
				sdi		=>	sdi,
				mode	=>	mode,
				hiz_b	=>	hiz_b,
				sdo		=>	sdo,
				dout1	=>	DIN1_zd,
				dout0	=>	DIN0_zd,
				ddr1	=>	DOUT1_ipd,
				ddr0	=>	DOUT0_ipd,
				padin	=>	padin,
				padout	=>	padout,
				padoen	=>	padoen,
				cbit	=>	pin_cbit
				);
				
	VITALTimingCheck : process (DOUT1_ipd,DOUT0_ipd,CLOCKENABLE_ipd,LATCHINPUTVALUE_ipd ,INPUTCLK_ipd ,OUTPUTENABLE_ipd, OUTPUTCLK_ipd,PACKAGEPIN_ipd , DIN1_zd,DIN0_zd ,PACKAGEPIN_zd )
			variable Tviol_CLOCKENABLE_INPUTCLK_posedge  :std_ulogic    := '0';
			variable Tviol_CLOCKENABLE_OUTPUTCLK_posedge  :std_ulogic    := '0';
			variable Tviol_PACKAGEPIN_INPUTCLK_posedge  :std_ulogic    := '0';
			variable Tviol_PACKAGEPIN_INPUTCLK_negedge  :std_ulogic    := '0';
			variable Tviol_PACKAGEPIN_OUTPUTCLK_posedge  :std_ulogic    := '0';
			variable Tviol_DOUT0_OUTPUTCLK_posedge  :std_ulogic    := '0';
			variable Tviol_DOUT0_OUTPUTCLK_negedge  :std_ulogic    := '0';
			variable Tviol_DOUT1_OUTPUTCLK_posedge  :std_ulogic    := '0';
			variable Tviol_DOUT1_OUTPUTCLK_negedge  :std_ulogic    := '0';
			variable Tviol_OUTPUTENABLE_OUTPUTCLK_posedge  :std_ulogic    := '0';
			
			variable Tmkr_CLOCKENABLE_INPUTCLK_posedge  :VitalTimingDataType    := VitalTimingDataInit;
			variable Tmkr_CLOCKENABLE_OUTPUTCLK_posedge  :VitalTimingDataType    := VitalTimingDataInit;
			variable Tmkr_PACKAGEPIN_INPUTCLK_posedge  :VitalTimingDataType    := VitalTimingDataInit;
			variable Tmkr_PACKAGEPIN_INPUTCLK_negedge  :VitalTimingDataType    := VitalTimingDataInit;
			variable Tmkr_PACKAGEPIN_OUTPUTCLK_posedge  :VitalTimingDataType    := VitalTimingDataInit;
			variable Tmkr_DOUT0_OUTPUTCLK_posedge  :VitalTimingDataType    := VitalTimingDataInit;
			variable Tmkr_DOUT0_OUTPUTCLK_negedge  :VitalTimingDataType    := VitalTimingDataInit;
			variable Tmkr_DOUT1_OUTPUTCLK_posedge  :VitalTimingDataType    := VitalTimingDataInit;
			variable Tmkr_DOUT1_OUTPUTCLK_negedge  :VitalTimingDataType    := VitalTimingDataInit;
			variable Tmkr_OUTPUTENABLE_OUTPUTCLK_posedge  :VitalTimingDataType    := VitalTimingDataInit;

begin
if (TimingChecksOn) then
			VitalSetupHoldCheck (
			Violation      => Tviol_CLOCKENABLE_INPUTCLK_posedge,
			TimingData     => Tmkr_CLOCKENABLE_INPUTCLK_posedge,
			TestSignal     => CLOCKENABLE_ipd,
			TestSignalName => "CLOCKENABLE",
			RefSignal      => INPUTCLK_ipd,
			RefSignalName  => "INPUTCLK",
			SetupHigh      => tsetup_CLOCKENABLE_INPUTCLK_posedge_posedge,
			SetupLow       => tsetup_CLOCKENABLE_INPUTCLK_negedge_posedge,
			HoldLow        => thold_CLOCKENABLE_INPUTCLK_posedge_posedge,
			HoldHigh       => thold_CLOCKENABLE_INPUTCLK_negedge_posedge,
			CheckEnabled   => true,
			RefTransition  => 'R',
			HeaderMsg      => "/SB_I0_OD",
			Xon            => Xon,
			MsgOn          => true,
			MsgSeverity    => warning);
			
				VitalSetupHoldCheck (
			Violation      => Tviol_CLOCKENABLE_OUTPUTCLK_posedge,
			TimingData     => Tmkr_CLOCKENABLE_OUTPUTCLK_posedge,
			TestSignal     => CLOCKENABLE_ipd,
			TestSignalName => "CLOCKENABLE",
			RefSignal      => OUTPUTCLK_ipd,
			RefSignalName  => "OUTPUTCLK",
			SetupHigh      => tsetup_CLOCKENABLE_OUTPUTCLK_posedge_posedge,
			SetupLow       => tsetup_CLOCKENABLE_OUTPUTCLK_negedge_posedge,
			HoldLow        => thold_CLOCKENABLE_OUTPUTCLK_posedge_posedge,
			HoldHigh       => thold_CLOCKENABLE_OUTPUTCLK_negedge_posedge,
			CheckEnabled   => true,
			RefTransition  => 'R',
			HeaderMsg      => "/SB_I0_OD",
			Xon            => Xon,
			MsgOn          => true,
			MsgSeverity    => warning);
			
			VitalSetupHoldCheck (
			Violation      => Tviol_OUTPUTENABLE_OUTPUTCLK_posedge,
			TimingData     => Tmkr_OUTPUTENABLE_OUTPUTCLK_posedge,
			TestSignal     => OUTPUTENABLE_ipd,
			TestSignalName => "OUTPUTENABLE",
			RefSignal      => OUTPUTCLK_ipd,
			RefSignalName  => "OUTPUTCLK",
			SetupHigh      => tsetup_OUTPUTENABLE_OUTPUTCLK_posedge_posedge,
			SetupLow       => tsetup_OUTPUTENABLE_OUTPUTCLK_negedge_posedge,
			HoldLow        => thold_OUTPUTENABLE_OUTPUTCLK_posedge_posedge,
			HoldHigh       => thold_OUTPUTENABLE_OUTPUTCLK_negedge_posedge,
			CheckEnabled   => true,
			RefTransition  => 'R',
			HeaderMsg      => "/SB_I0_OD",
			Xon            => Xon,
			MsgOn          => true,
			MsgSeverity    => warning);

	
	VitalSetupHoldCheck (
			Violation      => Tviol_PACKAGEPIN_INPUTCLK_posedge,
			TimingData     => Tmkr_PACKAGEPIN_INPUTCLK_posedge,
			TestSignal     => PACKAGEPIN_ipd,
			TestSignalName => "PACKAGEPIN",
			RefSignal      => INPUTCLK_ipd,
			RefSignalName  => "INPUTCLK",
			SetupHigh      => tsetup_PACKAGEPIN_INPUTCLK_posedge_posedge,
			SetupLow       => tsetup_PACKAGEPIN_INPUTCLK_negedge_posedge,
			HoldLow        => thold_PACKAGEPIN_INPUTCLK_posedge_posedge,
			HoldHigh       => thold_PACKAGEPIN_INPUTCLK_negedge_posedge,
			CheckEnabled   => true,
			RefTransition  => 'R',
			HeaderMsg      => "/SB_I0_OD",
			Xon            => Xon,
			MsgOn          => true,
			MsgSeverity    => warning);
			
			VitalSetupHoldCheck (
			Violation      => Tviol_PACKAGEPIN_INPUTCLK_negedge,
			TimingData     => Tmkr_PACKAGEPIN_INPUTCLK_negedge,
			TestSignal     => PACKAGEPIN_ipd,
			TestSignalName => "PACKAGEPIN",
			RefSignal      => INPUTCLK_ipd,
			RefSignalName  => "INPUTCLK",
			SetupHigh      => tsetup_PACKAGEPIN_INPUTCLK_posedge_negedge,
			SetupLow       => tsetup_PACKAGEPIN_INPUTCLK_negedge_negedge,
			HoldLow        => thold_PACKAGEPIN_INPUTCLK_posedge_negedge,
			HoldHigh       => thold_PACKAGEPIN_INPUTCLK_negedge_negedge,
			CheckEnabled   => true,
			RefTransition  => 'F',
			HeaderMsg      => "/SB_I0_OD",
			Xon            => Xon,
			MsgOn          => true,
			MsgSeverity    => warning);
			
				VitalSetupHoldCheck (
			Violation      => Tviol_PACKAGEPIN_INPUTCLK_negedge,
			TimingData     => Tmkr_PACKAGEPIN_INPUTCLK_negedge,
			TestSignal     => PACKAGEPIN_ipd,
			TestSignalName => "PACKAGEPIN",
			RefSignal      => INPUTCLK_ipd,
			RefSignalName  => "INPUTCLK",
			SetupHigh      => tsetup_PACKAGEPIN_INPUTCLK_posedge_negedge,
			SetupLow       => tsetup_PACKAGEPIN_INPUTCLK_negedge_negedge,
			HoldLow        => thold_PACKAGEPIN_INPUTCLK_posedge_negedge,
			HoldHigh       => thold_PACKAGEPIN_INPUTCLK_negedge_negedge,
			CheckEnabled   => true,
			RefTransition  => 'F',
			HeaderMsg      => "/SB_I0_OD",
			Xon            => Xon,
			MsgOn          => true,
			MsgSeverity    => warning);
			
			
			VitalSetupHoldCheck (
			Violation      => Tviol_PACKAGEPIN_OUTPUTCLK_posedge,
			TimingData     => Tmkr_PACKAGEPIN_OUTPUTCLK_posedge,
			TestSignal     => PACKAGEPIN_ipd,
			TestSignalName => "PACKAGEPIN",
			RefSignal      => OUTPUTCLK_ipd,
			RefSignalName  => "OUTPUTCLK",
			SetupHigh      => tsetup_PACKAGEPIN_OUTPUTCLK_posedge_posedge,
			SetupLow       => tsetup_PACKAGEPIN_OUTPUTCLK_negedge_posedge,
			HoldLow        => thold_PACKAGEPIN_OUTPUTCLK_posedge_posedge,
			HoldHigh       => thold_PACKAGEPIN_OUTPUTCLK_negedge_posedge,
			CheckEnabled   => true,
			RefTransition  => 'R',
			HeaderMsg      => "/SB_I0_OD",
			Xon            => Xon,
			MsgOn          => true,
			MsgSeverity    => warning);
			
			
				VitalSetupHoldCheck (
			Violation      => Tviol_DOUT0_OUTPUTCLK_posedge,
			TimingData     => Tmkr_DOUT0_OUTPUTCLK_posedge,
			TestSignal     => DOUT0_ipd,
			TestSignalName => "DOUT0",
			RefSignal      => OUTPUTCLK_ipd,
			RefSignalName  => "OUTPUTCLK",
			SetupHigh      => tsetup_DOUT0_OUTPUTCLK_posedge_posedge,
			SetupLow       => tsetup_DOUT0_OUTPUTCLK_negedge_posedge,
			HoldLow        => thold_DOUT0_OUTPUTCLK_posedge_posedge,
			HoldHigh       => thold_DOUT0_OUTPUTCLK_negedge_posedge,
			CheckEnabled   => true,
			RefTransition  => 'R',
			HeaderMsg      => "/SB_I0_OD",
			Xon            => Xon,
			MsgOn          => true,
			MsgSeverity    => warning);
			
			
			VitalSetupHoldCheck (
			Violation      => Tviol_DOUT1_OUTPUTCLK_posedge,
			TimingData     => Tmkr_DOUT1_OUTPUTCLK_posedge,
			TestSignal     => DOUT1_ipd,
			TestSignalName => "DOUT1",
			RefSignal      => OUTPUTCLK_ipd,
			RefSignalName  => "OUTPUTCLK",
			SetupHigh      => tsetup_DOUT1_OUTPUTCLK_posedge_posedge,
			SetupLow       => tsetup_DOUT1_OUTPUTCLK_negedge_posedge,
			HoldLow        => thold_DOUT1_OUTPUTCLK_posedge_posedge,
			HoldHigh       => thold_DOUT1_OUTPUTCLK_negedge_posedge,
			CheckEnabled   => true,
			RefTransition  => 'R',
			HeaderMsg      => "/SB_I0_OD",
			Xon            => Xon,
			MsgOn          => true,
			MsgSeverity    => warning);
			
			VitalSetupHoldCheck (
			Violation      => Tviol_DOUT1_OUTPUTCLK_negedge,
			TimingData     => Tmkr_DOUT1_OUTPUTCLK_negedge,
			TestSignal     => DOUT1_ipd,
			TestSignalName => "DOUT1",
			RefSignal      => OUTPUTCLK_ipd,
			RefSignalName  => "OUTPUTCLK",
			SetupHigh      => tsetup_DOUT1_OUTPUTCLK_posedge_negedge,
			SetupLow       => tsetup_DOUT1_OUTPUTCLK_negedge_negedge,
			HoldLow        => thold_DOUT1_OUTPUTCLK_posedge_negedge,
			HoldHigh       => thold_DOUT1_OUTPUTCLK_negedge_negedge,
			CheckEnabled   => true,
			RefTransition  => 'F',
			HeaderMsg      => "/SB_I0_OD",
			Xon            => Xon,
			MsgOn          => true,
			MsgSeverity    => warning);
			end if;
end process;
				
	VITALPathDelay :process (DOUT1_ipd,DOUT0_ipd,CLOCKENABLE_ipd,LATCHINPUTVALUE_ipd ,INPUTCLK_ipd ,OUTPUTENABLE_ipd, OUTPUTCLK_ipd,PACKAGEPIN_ipd , DIN1_zd,DIN0_zd ,PACKAGEPIN_zd )
	
	variable DIN0_GlitchData : VitalGlitchDataType;
	variable DIN1_GlitchData : VitalGlitchDataType;
	variable PACKAGEPIN_GlitchData : VitalGlitchDataType;
	variable DIN0_tmp : std_ulogic :='X';
	variable DIN1_tmp : std_ulogic :='X';
	variable PACKAGEPIN_tmp : std_ulogic :='X';
	begin	  
		DIN0_tmp:=DIN0_zd;
		DIN1_tmp:=DIN1_zd; 
		PACKAGEPIN_tmp:=PACKAGEPIN_zd;
VitalPathDelay01 (
      OutSignal                 => DIN0,
      GlitchData                => DIN0_GlitchData,
      OutSignalName             => "DIN0",
      OutTemp                   => DIN0_tmp,
      Paths                     => (0 =>(PACKAGEPIN_ipd'last_event, tpd_PACKAGEPIN_DIN0, true),
									1 =>(LATCHINPUTVALUE_ipd'last_event, tpd_LATCHINPUTVALUE_DIN0, true),
									2 =>(INPUTCLK_ipd'last_event, tpd_INPUTCLK_DIN0_posedge, true)),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
VitalPathDelay01 (
      OutSignal                 => DIN1,
      GlitchData                => DIN1_GlitchData,
      OutSignalName             => "DIN1",
      OutTemp                   => DIN1_tmp,
      Paths                     => (0 =>(PACKAGEPIN_ipd'last_event, tpd_PACKAGEPIN_DIN1, true),
									1 =>(LATCHINPUTVALUE_ipd'last_event, tpd_LATCHINPUTVALUE_DIN1, true),
									2 =>(INPUTCLK_ipd'last_event, tpd_INPUTCLK_DIN1_negedge, true)),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
VitalPathDelay01 (
      OutSignal                 => PACKAGEPIN,
      GlitchData                => PACKAGEPIN_GlitchData,
      OutSignalName             => "PACKAGEPIN",
      OutTemp                   => PACKAGEPIN_tmp,
      Paths                     => (0 =>(DOUT0_ipd'last_event, tpd_DOUT0_PACKAGEPIN, true),
									1 =>(DOUT1_ipd'last_event, tpd_DOUT1_PACKAGEPIN, true),
									2 =>(OUTPUTENABLE_ipd'last_event, tpd_OUTPUTENABLE_PACKAGEPIN, true),
									3 =>(OUTPUTCLK_ipd'last_event, tpd_OUTPUTCLK_PACKAGEPIN, true),
									4 =>(INPUTCLK_ipd'last_event, tpd_INPUTCLK_PACKAGEPIN, true)),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);

end process;

end	SB_IO_OD_V;

-----------------------------------------------------
---     	SB_HFOSC 		-------
------------------------------------------------
library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use IEEE.Vital_Primitives.all;
use IEEE.VITAL_Timing.all;
entity  SB_HFOSC  is 
	generic( CLKHF_DIV: string:="0b00";
				Xon   : boolean := true;
				MsgOn : boolean := true;
				tipd_CLKHFEN: VitalDelayType01 := (0.000 ns, 0.000 ns);
				tipd_CLKHFPU: VitalDelayType01 := (0.000 ns, 0.000 ns);
				tpd_CLKHFEN_CLKHF : VitalDelayType01 := (0.000 ns, 0.000 ns);
				tpd_CLKHFPU_CLKHF : VitalDelayType01 := (0.000 ns, 0.000 ns)
); 
port(
	CLKHF : out std_logic;
	CLKHFEN  :in std_logic;
    CLKHFPU : in std_logic
    );
		attribute VITAL_LEVEL0 of			    
    SB_HFOSC  : entity is true;
end SB_HFOSC ;

architecture SB_HFOSC_V of SB_HFOSC is
attribute VITAL_LEVEL0 of
    SB_HFOSC_V : architecture is true;
	signal CLKHFEN_ipd: std_ulogic := 'X';
	signal CLKHFPU_ipd: std_ulogic := 'X';
	signal CLKHF_sig  : std_ulogic	:='X';
  
component SB_HFOSC_CORE				    
generic( CLKHF_DIV: string:="0b00"); 	
port ( 
	CLKHF_PU : IN std_logic;
	CLKHF_EN : IN std_logic;
	CLKHF : OUT std_logic
);

end component;

begin
WireDelay : block
  begin
    VitalWireDelay (CLKHFEN_ipd, CLKHFEN, tipd_CLKHFEN);
	VitalWireDelay (CLKHFPU_ipd, CLKHFPU, tipd_CLKHFPU);
  end block;

LS: SB_HFOSC_CORE 					 
GENERIC MAP (CLKHF_DIV => CLKHF_DIV)
port map(
	CLKHF_PU=> CLKHFPU_ipd,
	CLKHF_EN=> CLKHFEN,
	CLKHF=> CLKHF_sig
		);
VITALPathDelay :process (CLKHFEN_ipd,CLKHF_sig,CLKHFPU_ipd)
variable CLKHF_GlitchData : VitalGlitchDataType;  
variable CLKHF_zd  : std_ulogic	:='X';
begin  
	CLKHF_zd:=CLKHF_sig;
VitalPathDelay01 (
      OutSignal                 => CLKHF,
      GlitchData                => CLKHF_GlitchData,
      OutSignalName             => "CLKHF",
      OutTemp                   => CLKHF_zd,
      Paths                     => (--0 =>(CLKHFEN_ipd'last_event, tpd_CLKHFEN_CLKHF, true),
									0 =>(CLKHFPU_ipd'last_event, tpd_CLKHFPU_CLKHF, true)),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
end process;

end 	SB_HFOSC_V; 

--------------------------------------------------------------
---     	SB_LFOSC 		-------
------------------------------------------------

library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use IEEE.Vital_Primitives.all;
use IEEE.VITAL_Timing.all;
entity  SB_LFOSC  is 
generic(
	Xon   : boolean := true;
    MsgOn : boolean := true;
	tipd_CLKLFEN: VitalDelayType01 := (0.000 ns, 0.000 ns);
	tipd_CLKLFPU: VitalDelayType01 := (0.000 ns, 0.000 ns);
	tpd_CLKLFEN_CLKLF : VitalDelayType01 := (0.000 ns, 0.000 ns);
    tpd_CLKLFPU_CLKLF : VitalDelayType01 := (0.000 ns, 0.000 ns)
 ); 
port(
	CLKLF : out std_logic;
	CLKLFEN  :in std_logic;
    CLKLFPU : in std_logic
    );
	attribute VITAL_LEVEL0 of			    
    SB_LFOSC  : entity is true;
end SB_LFOSC ;

architecture SB_LFOSC_V of SB_LFOSC is
attribute VITAL_LEVEL0 of
    SB_LFOSC_V : architecture is true;
	signal CLKLFEN_ipd: std_ulogic := 'X';
	signal CLKLFPU_ipd: std_ulogic := 'X';
	signal CLKLF_sig  : std_ulogic	:='X';
  
component SB_LFOSC_CORE		
port ( 
	CLKLF_PU : IN std_logic;
	CLKLF_EN : IN std_logic;
	CLKLF : OUT std_logic
);
end component;

begin

WireDelay : block
  begin
    VitalWireDelay (CLKLFEN_ipd, CLKLFEN, tipd_CLKLFEN);
	VitalWireDelay (CLKLFPU_ipd, CLKLFPU, tipd_CLKLFPU);
  end block;

LS: SB_LFOSC_CORE 
port map(
	CLKLF_PU=> CLKLFPU_ipd,
	CLKLF_EN=> CLKLFEN,
	CLKLF=> CLKLF_sig
		);
		
VITALPathDelay :process (CLKLFEN_ipd,CLKLF_sig,CLKLFPU_ipd)
variable CLKLF_GlitchData : VitalGlitchDataType;
variable CLKLF_zd  : std_ulogic	:='X';
begin		  
	CLKLF_zd:=CLKLF_sig;
VitalPathDelay01 (
      OutSignal                 => CLKLF,
      GlitchData                => CLKLF_GlitchData,
      OutSignalName             => "CLKLF",
      OutTemp                   => CLKLF_zd,
      Paths                     => (--0 =>(CLKLFEN_ipd'last_event, tpd_CLKLFEN_CLKLF, true),
									0 =>(CLKLFPU_ipd'last_event, tpd_CLKLFPU_CLKLF, true)),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
end process;

end 	SB_LFOSC_V; 


-------------------------------------------------
---     	SB_IR_DRV 		-------
------------------------------------------------

library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;
entity  SB_IR_DRV  is 
	generic( 
		TimingChecksOn : boolean := true;
        Xon            : boolean := false;
        MsgOn          : boolean := false;
		tipd_IRLEDEN: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_IRPU: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_IRPWM: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tpd_IRPWM_IRLED : VitalDelayType01 := (0.000 ns, 0.000 ns);
		IR_CURRENT: string:="0b0000000000" ); 
port(
	IRLED : out std_logic;
	IRLEDEN  :in std_logic;
	IRPU  :in std_logic;						 
    IRPWM : in std_logic
    );
	attribute VITAL_LEVEL0 of			    
    SB_IR_DRV  : entity is true;
end SB_IR_DRV ;

architecture SB_IR_DRV_V of SB_IR_DRV is
attribute VITAL_LEVEL0 of
    SB_IR_DRV_V : architecture is true; 
	signal IRPU_ipd: std_ulogic := 'X';
	signal IRLEDEN_ipd: std_ulogic := 'X';
	signal IRPWM_ipd: std_ulogic := 'X';
	signal IRLED_sig  : std_ulogic	:='X';
component  SB_IR_DRV_CORE
	generic( IR_CURRENT: string:="0b0000000000" ); 
port(
	IRLED : out std_logic;
	IRLED_EN  :in std_logic;
	IR_PU  :in std_logic;
    IR_PWM : in std_logic
    );
end component;

begin
WireDelay : block
  begin
    VitalWireDelay (IRLEDEN_ipd, IRLEDEN, tipd_IRLEDEN);
	VitalWireDelay (IRPU_ipd, IRPU, tipd_IRPU);
	VitalWireDelay (IRPWM_ipd, IRPWM, tipd_IRPWM);
  end block;
LS: SB_IR_DRV_CORE 
generic map( IR_CURRENT=>IR_CURRENT )
port map(
	IRLED =>IRLED_sig,
	IRLED_EN=>IRLEDEN_ipd,  
	IR_PU=>IRPU_ipd,  
    IR_PWM=> IRPWM_ipd 
);
VITALPathDelay :process (IRPWM_ipd,IRPU_ipd,IRLEDEN_ipd,IRLED_sig)
variable IRLED_GlitchData : VitalGlitchDataType; 
variable IRLED_zd : std_ulogic :='X';
begin										  
	IRLED_zd:=IRLED_sig;
VitalPathDelay01 (
      OutSignal                 => IRLED,
      GlitchData                => IRLED_GlitchData,
      OutSignalName             => "IRLED",
      OutTemp                   => IRLED_zd,
      Paths                     => (0 =>(IRPWM_ipd'last_event, tpd_IRPWM_IRLED, true)),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
end process;
end 	SB_IR_DRV_V; 

--------------------------------------------------
---     	SB_LEDD_IP 		-------
------------------------------------------------

library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;
entity  SB_LEDD_IP  is 

generic (
	TimingChecksOn  	: boolean := true;
	Xon   			: boolean := true;
	MsgOn 			: boolean := true;

	tipd_LEDDCS:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDCLK:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDDAT7:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDDAT6:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDDAT5:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDDAT4:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDDAT3:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDDAT2:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDDAT1:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDDAT0:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDADDR3:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDADDR2:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDADDR1:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDADDR0:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDDEN:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDEXE:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDRST:VitalDelayType01 := (0 ns, 0 ns);
	tpd_LEDDCLK_LEDDON_posedge :VitalDelayType01 := (100 ns, 100 ns);
	tpd_LEDDCLK_PWMOUT0_posedge :VitalDelayType01 := (100 ns, 100 ns);
	tpd_LEDDCLK_PWMOUT1_posedge :VitalDelayType01 := (100 ns, 100 ns);
	tpd_LEDDCLK_PWMOUT2_posedge :VitalDelayType01 := (100 ns, 100 ns);
	
	tsetup_LEDDCS_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;	
	tsetup_LEDDCS_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDEN_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;	
	tsetup_LEDDDEN_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDEXE_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;	
	tsetup_LEDDEXE_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDADDR0_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDADDR0_LEDDCLK_negedge_posedge :VitalDelayType := 0 ns;
	tsetup_LEDDADDR1_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDADDR1_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDADDR2_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDADDR2_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDADDR3_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDADDR3_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	
	tsetup_LEDDDAT0_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDAT0_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDAT1_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDAT1_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDAT2_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDAT2_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDAT3_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDAT3_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDAT4_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDAT4_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDAT5_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDAT5_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDAT6_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDAT6_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDAT7_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDAT7_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	
	thold_LEDDCS_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;	
	thold_LEDDCS_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDEN_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;	
	thold_LEDDDEN_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDEXE_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;	
	thold_LEDDEXE_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDADDR0_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDADDR0_LEDDCLK_negedge_posedge :VitalDelayType := 0 ns;
	thold_LEDDADDR1_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDADDR1_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDADDR2_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDADDR2_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDADDR3_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDADDR3_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	
	thold_LEDDDAT0_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDAT0_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDAT1_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDAT1_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDAT2_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDAT2_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDAT3_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDAT3_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDAT4_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDAT4_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDAT5_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDAT5_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDAT6_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDAT6_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDAT7_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDAT7_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns
	
);
 
port(
	PWMOUT0 : out std_logic;	
	PWMOUT1 : out std_logic;
	PWMOUT2 : out std_logic;
	LEDDON : out std_logic; 
	LEDDCS:in std_logic;
	LEDDCLK:in std_logic;
	LEDDDAT7:in std_logic;
	LEDDDAT6:in std_logic;
	LEDDDAT5:in std_logic;
	LEDDDAT4:in std_logic;
	LEDDDAT3:in std_logic;
	LEDDDAT2:in std_logic;
	LEDDDAT1:in std_logic;
	LEDDDAT0:in std_logic;
	LEDDADDR3:in std_logic;
	LEDDADDR2:in std_logic;
	LEDDADDR1:in std_logic;
	LEDDADDR0:in std_logic;
	LEDDDEN:in std_logic;
	LEDDEXE:in std_logic;
	LEDDRST:in std_logic
    );
	attribute VITAL_LEVEL0 of			    
    SB_LEDD_IP  : entity is true;
end SB_LEDD_IP ;

architecture SB_LEDD_IP_V of SB_LEDD_IP is
attribute VITAL_LEVEL0 of
    SB_LEDD_IP_V : architecture is true;

SIGNAL LEDD_ADDR: std_logic_vector (3 downto 0);   
SIGNAL LEDD_DAT: std_logic_vector (7 downto 0);

	signal  PWMOUT0_sig  : std_ulogic	:='X';	
	signal  PWMOUT1_sig  : std_ulogic	:='X';
	signal  PWMOUT2_sig  : std_ulogic	:='X';
	signal  LEDDON_sig  : std_ulogic	:='X'; 
	
	signal  LEDDCS_ipd: std_ulogic := 'X';
	signal  LEDDCLK_ipd: std_ulogic := 'X';
	signal  LEDDDAT7_ipd: std_ulogic := 'X';
	signal  LEDDDAT6_ipd: std_ulogic := 'X';
	signal  LEDDDAT5_ipd: std_ulogic := 'X';
	signal  LEDDDAT4_ipd: std_ulogic := 'X';
	signal  LEDDDAT3_ipd: std_ulogic := 'X';
	signal  LEDDDAT2_ipd: std_ulogic := 'X';
	signal  LEDDDAT1_ipd: std_ulogic := 'X';
	signal  LEDDDAT0_ipd: std_ulogic := 'X';
	signal  LEDDADDR3_ipd: std_ulogic := 'X';
	signal  LEDDADDR2_ipd: std_ulogic := 'X';
	signal  LEDDADDR1_ipd: std_ulogic := 'X';
	signal  LEDDADDR0_ipd: std_ulogic := 'X';
	signal  LEDDDEN_ipd: std_ulogic := 'X';
	signal  LEDDEXE_ipd: std_ulogic := 'X';
	signal  LEDDRST_ipd: std_ulogic := 'X';
    	signal  ledd_rst   : std_logic := '1';
component ledd_ip 
port	(
	pwm_out_r:out std_logic;
	pwm_out_g:out std_logic;
	pwm_out_b:out std_logic; 
	ledd_on :out std_logic;
	ledd_rst_async :in std_logic; 
	ledd_clk :in std_logic;
	ledd_cs :in std_logic;
	ledd_den :in std_logic; 
	ledd_adr :in std_logic_vector (3 downto 0); 
	ledd_dat :in std_logic_vector (7 downto 0);
    ledd_exe :in std_logic
   );
end component;

begin
	-- device reset of irip for 100ns --- 
process 
    begin
            wait for 100 ns;
            ledd_rst <= '0';
	    wait; 
end process;


WireDelay : block
  begin
    VitalWireDelay (LEDDCS_ipd, LEDDCS, tipd_LEDDCS);
	VitalWireDelay (LEDDCLK_ipd, LEDDCLK, tipd_LEDDCLK);
	VitalWireDelay (LEDDDAT7_ipd, LEDDDAT7, tipd_LEDDDAT7);
	VitalWireDelay (LEDDDAT6_ipd, LEDDDAT6, tipd_LEDDDAT6);
	VitalWireDelay (LEDDDAT5_ipd, LEDDDAT5, tipd_LEDDDAT5);
	VitalWireDelay (LEDDDAT4_ipd, LEDDDAT4, tipd_LEDDDAT4);
	VitalWireDelay (LEDDDAT3_ipd, LEDDDAT3, tipd_LEDDDAT3);
	VitalWireDelay (LEDDDAT2_ipd, LEDDDAT2, tipd_LEDDDAT2);
	VitalWireDelay (LEDDDAT1_ipd, LEDDDAT1, tipd_LEDDDAT1);
	VitalWireDelay (LEDDDAT0_ipd, LEDDDAT0, tipd_LEDDDAT0);
	VitalWireDelay (LEDDADDR3_ipd, LEDDADDR3, tipd_LEDDADDR3);
	VitalWireDelay (LEDDADDR2_ipd, LEDDADDR2, tipd_LEDDADDR2);
	VitalWireDelay (LEDDADDR1_ipd, LEDDADDR1, tipd_LEDDADDR1);
	VitalWireDelay (LEDDADDR0_ipd, LEDDADDR0, tipd_LEDDADDR0);
	VitalWireDelay (LEDDDEN_ipd, LEDDDEN, tipd_LEDDDEN);
	VitalWireDelay (LEDDEXE_ipd, LEDDEXE, tipd_LEDDEXE);
	VitalWireDelay (LEDDRST_ipd, LEDDRST, tipd_LEDDRST);
	
  end block;

LS: ledd_ip 
port map(
	pwm_out_r =>PWMOUT0_sig  ,
	pwm_out_g =>PWMOUT1_sig  ,
	pwm_out_b =>PWMOUT2_sig  , 
	ledd_on  =>LEDDON_sig  ,
	ledd_rst_async  =>ledd_rst  , 
	ledd_clk  => LEDDCLK_ipd ,
	ledd_cs  => LEDDCS_ipd ,
	ledd_den  => LEDDDEN_ipd , 
	ledd_adr =>LEDD_ADDR,    
	ledd_dat  =>LEDD_DAT,    
    ledd_exe => LEDDEXE_ipd   
);
LEDD_ADDR<=(LEDDADDR3_ipd,LEDDADDR2_ipd,LEDDADDR1_ipd,LEDDADDR0_ipd) ; 
LEDD_DAT<=(LEDDDAT7_ipd,LEDDDAT6_ipd,LEDDDAT5_ipd,LEDDDAT4_ipd,LEDDDAT3_ipd,LEDDDAT2_ipd,LEDDDAT1_ipd,LEDDDAT0_ipd);

VITALBehavior : process(  PWMOUT0_sig,PWMOUT1_sig, PWMOUT2_sig,LEDDON_sig,LEDDCS_ipd,LEDDCLK_ipd,LEDDDAT7_ipd,LEDDDAT6_ipd,
	  LEDDDAT5_ipd,LEDDDAT4_ipd,LEDDDAT3_ipd,LEDDDAT2_ipd,LEDDDAT1_ipd,LEDDDAT0_ipd,LEDDADDR3_ipd,LEDDADDR2_ipd,LEDDADDR1_ipd,
	  LEDDADDR0_ipd,LEDDDEN_ipd,LEDDEXE_ipd,LEDDRST_ipd)

	variable Tviol_LEDDCS_LEDDCLK_posedge : std_logic := '0';	
	variable Tviol_LEDDDEN_LEDDCLK_posedge : std_logic := '0';	
	variable Tviol_LEDDEXE_LEDDCLK_posedge : std_logic := '0';	
	variable Tviol_LEDDADDR0_LEDDCLK_posedge : std_logic := '0';
	variable Tviol_LEDDADDR1_LEDDCLK_posedge : std_logic := '0';
	variable Tviol_LEDDADDR2_LEDDCLK_posedge : std_logic := '0';
	variable Tviol_LEDDADDR3_LEDDCLK_posedge : std_logic := '0';

	variable Tviol_LEDDDAT0_LEDDCLK_posedge : std_logic := '0';
	variable Tviol_LEDDDAT1_LEDDCLK_posedge : std_logic := '0';
	variable Tviol_LEDDDAT2_LEDDCLK_posedge : std_logic := '0';
	variable Tviol_LEDDDAT3_LEDDCLK_posedge : std_logic := '0';
	variable Tviol_LEDDDAT4_LEDDCLK_posedge : std_logic := '0';
	variable Tviol_LEDDDAT5_LEDDCLK_posedge : std_logic := '0';
	variable Tviol_LEDDDAT6_LEDDCLK_posedge : std_logic := '0';
	variable Tviol_LEDDDAT7_LEDDCLK_posedge : std_logic := '0';
	
	variable Tmkr_LEDDCS_LEDDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;	
	variable Tmkr_LEDDDEN_LEDDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;	
	variable Tmkr_LEDDEXE_LEDDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;	
	variable Tmkr_LEDDADDR0_LEDDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LEDDADDR1_LEDDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LEDDADDR2_LEDDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LEDDADDR3_LEDDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;

	variable Tmkr_LEDDDAT0_LEDDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LEDDDAT1_LEDDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LEDDDAT2_LEDDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LEDDDAT3_LEDDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LEDDDAT4_LEDDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LEDDDAT5_LEDDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LEDDDAT6_LEDDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LEDDDAT7_LEDDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable LEDDON_GlitchData : VitalGlitchDataType;  
	variable PWMOUT0_GlitchData : VitalGlitchDataType;
	variable PWMOUT1_GlitchData : VitalGlitchDataType;
	variable PWMOUT2_GlitchData : VitalGlitchDataType;				 
	variable PWMOUT0_zd :std_ulogic :='X';
	variable PWMOUT1_zd :std_ulogic :='X';
	variable PWMOUT2_zd :std_ulogic :='X'; 
	variable LEDDON_zd : std_ulogic :='X';

begin	  	
	PWMOUT0_zd:=PWMOUT0_sig;
	PWMOUT1_zd:=PWMOUT1_sig;
	PWMOUT2_zd:=PWMOUT2_sig;
	LEDDON_zd :=LEDDON_sig;
	if (TimingChecksOn) then
      VitalSetupHoldCheck (
        Violation      => Tviol_LEDDCS_LEDDCLK_posedge,
        TimingData     => Tmkr_LEDDCS_LEDDCLK_posedge,
        TestSignal     => LEDDCS_ipd,
        TestSignalName => "LEDDCS",
        TestDelay      => 0 ns,
        RefSignal      => LEDDCLK_ipd,
        RefSignalName  => "LEDDCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_LEDDCS_LEDDCLK_posedge_posedge,
        SetupLow       => tsetup_LEDDCS_LEDDCLK_negedge_posedge,
        HoldLow        => thold_LEDDCS_LEDDCLK_posedge_posedge,
        HoldHigh       => thold_LEDDCS_LEDDCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_LEDD_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	  
	      VitalSetupHoldCheck (
        Violation      => Tviol_LEDDDEN_LEDDCLK_posedge,
        TimingData     => Tmkr_LEDDDEN_LEDDCLK_posedge,
        TestSignal     => LEDDDEN_ipd,
        TestSignalName => "LEDDDEN",
        TestDelay      => 0 ns,
        RefSignal      => LEDDCLK_ipd,
        RefSignalName  => "LEDDCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_LEDDDEN_LEDDCLK_posedge_posedge,
        SetupLow       => tsetup_LEDDDEN_LEDDCLK_negedge_posedge,
        HoldLow        => thold_LEDDDEN_LEDDCLK_posedge_posedge,
        HoldHigh       => thold_LEDDDEN_LEDDCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_LEDD_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	 
		
		      VitalSetupHoldCheck (
        Violation      => Tviol_LEDDEXE_LEDDCLK_posedge,
        TimingData     => Tmkr_LEDDEXE_LEDDCLK_posedge,
        TestSignal     => LEDDEXE_ipd,
        TestSignalName => "LEDDEXE",
        TestDelay      => 0 ns,
        RefSignal      => LEDDCLK_ipd,
        RefSignalName  => "LEDDCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_LEDDEXE_LEDDCLK_posedge_posedge,
        SetupLow       => tsetup_LEDDEXE_LEDDCLK_negedge_posedge,
        HoldLow        => thold_LEDDEXE_LEDDCLK_posedge_posedge,
        HoldHigh       => thold_LEDDEXE_LEDDCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_LEDD_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	 
		
		      VitalSetupHoldCheck (
        Violation      => Tviol_LEDDADDR0_LEDDCLK_posedge,
        TimingData     => Tmkr_LEDDADDR0_LEDDCLK_posedge,
        TestSignal     => LEDDADDR0_ipd,	 
        TestSignalName => "LEDDADDR0",
        TestDelay      => 0 ns,
        RefSignal      => LEDDCLK_ipd,
        RefSignalName  => "LEDDCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_LEDDADDR0_LEDDCLK_posedge_posedge,
        SetupLow       => tsetup_LEDDADDR0_LEDDCLK_negedge_posedge,
        HoldLow        => thold_LEDDADDR0_LEDDCLK_posedge_posedge,
        HoldHigh       => thold_LEDDADDR0_LEDDCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_LEDD_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	 
		
		      VitalSetupHoldCheck (
        Violation      => Tviol_LEDDADDR1_LEDDCLK_posedge,
        TimingData     => Tmkr_LEDDADDR1_LEDDCLK_posedge,
        TestSignal     => LEDDADDR1_ipd,
        TestSignalName => "LEDDADDR1",
        TestDelay      => 0 ns,
        RefSignal      => LEDDCLK_ipd,
        RefSignalName  => "LEDDCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_LEDDADDR1_LEDDCLK_posedge_posedge,
        SetupLow       => tsetup_LEDDADDR1_LEDDCLK_negedge_posedge,
        HoldLow        => thold_LEDDADDR1_LEDDCLK_posedge_posedge,
        HoldHigh       => thold_LEDDADDR1_LEDDCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_LEDD_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
		
		      VitalSetupHoldCheck (
        Violation      => Tviol_LEDDADDR2_LEDDCLK_posedge,
        TimingData     => Tmkr_LEDDADDR2_LEDDCLK_posedge,
        TestSignal     => LEDDADDR2_ipd,
        TestSignalName => "LEDDADDR2",
        TestDelay      => 0 ns,
        RefSignal      => LEDDCLK_ipd,
        RefSignalName  => "LEDDCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_LEDDADDR2_LEDDCLK_posedge_posedge,
        SetupLow       => tsetup_LEDDADDR2_LEDDCLK_negedge_posedge,
        HoldLow        => thold_LEDDADDR2_LEDDCLK_posedge_posedge,
        HoldHigh       => thold_LEDDADDR2_LEDDCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_LEDD_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
		
		      VitalSetupHoldCheck (
        Violation      => Tviol_LEDDADDR3_LEDDCLK_posedge,
        TimingData     => Tmkr_LEDDADDR3_LEDDCLK_posedge,
        TestSignal     => LEDDADDR3_ipd,
        TestSignalName => "LEDDADDR3",
        TestDelay      => 0 ns,
        RefSignal      => LEDDCLK_ipd,
        RefSignalName  => "LEDDCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_LEDDADDR3_LEDDCLK_posedge_posedge,
        SetupLow       => tsetup_LEDDADDR3_LEDDCLK_negedge_posedge,
        HoldLow        => thold_LEDDADDR3_LEDDCLK_posedge_posedge,
        HoldHigh       => thold_LEDDADDR3_LEDDCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_LEDD_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);		 
		
		   VitalSetupHoldCheck (
        Violation      => Tviol_LEDDDAT0_LEDDCLK_posedge,
        TimingData     => Tmkr_LEDDDAT0_LEDDCLK_posedge,
        TestSignal     => LEDDDAT0_ipd,
        TestSignalName => "LEDDDAT0",
        TestDelay      => 0 ns,
        RefSignal      => LEDDCLK_ipd,
        RefSignalName  => "LEDDCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_LEDDDAT0_LEDDCLK_posedge_posedge,
        SetupLow       => tsetup_LEDDDAT0_LEDDCLK_negedge_posedge,
        HoldLow        => thold_LEDDDAT0_LEDDCLK_posedge_posedge,
        HoldHigh       => thold_LEDDDAT0_LEDDCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_LEDD_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
		
		   VitalSetupHoldCheck (
        Violation      => Tviol_LEDDDAT1_LEDDCLK_posedge,
        TimingData     => Tmkr_LEDDDAT1_LEDDCLK_posedge,
        TestSignal     => LEDDDAT1_ipd,
        TestSignalName => "LEDDDAT1",
        TestDelay      => 0 ns,
        RefSignal      => LEDDCLK_ipd,
        RefSignalName  => "LEDDCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_LEDDDAT1_LEDDCLK_posedge_posedge,
        SetupLow       => tsetup_LEDDDAT1_LEDDCLK_negedge_posedge,
        HoldLow        => thold_LEDDDAT1_LEDDCLK_posedge_posedge,
        HoldHigh       => thold_LEDDDAT1_LEDDCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_LEDD_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
		
		   VitalSetupHoldCheck (
        Violation      => Tviol_LEDDDAT2_LEDDCLK_posedge,
        TimingData     => Tmkr_LEDDDAT2_LEDDCLK_posedge,
        TestSignal     => LEDDDAT2_ipd,
        TestSignalName => "LEDDDAT2",
        TestDelay      => 0 ns,
        RefSignal      => LEDDCLK_ipd,
        RefSignalName  => "LEDDCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_LEDDDAT2_LEDDCLK_posedge_posedge,
        SetupLow       => tsetup_LEDDDAT2_LEDDCLK_negedge_posedge,
        HoldLow        => thold_LEDDDAT2_LEDDCLK_posedge_posedge,
        HoldHigh       => thold_LEDDDAT2_LEDDCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_LEDD_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
		
		
		   VitalSetupHoldCheck (
        Violation      => Tviol_LEDDDAT3_LEDDCLK_posedge,
        TimingData     => Tmkr_LEDDDAT3_LEDDCLK_posedge,
        TestSignal     => LEDDDAT3_ipd,
        TestSignalName => "LEDDDAT3",
        TestDelay      => 0 ns,
        RefSignal      => LEDDCLK_ipd,
        RefSignalName  => "LEDDCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_LEDDDAT3_LEDDCLK_posedge_posedge,
        SetupLow       => tsetup_LEDDDAT3_LEDDCLK_negedge_posedge,
        HoldLow        => thold_LEDDDAT3_LEDDCLK_posedge_posedge,
        HoldHigh       => thold_LEDDDAT3_LEDDCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_LEDD_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
		
		
		   VitalSetupHoldCheck (
        Violation      => Tviol_LEDDDAT4_LEDDCLK_posedge,
        TimingData     => Tmkr_LEDDDAT4_LEDDCLK_posedge,
        TestSignal     => LEDDDAT4_ipd,
        TestSignalName => "LEDDDAT4",
        TestDelay      => 0 ns,
        RefSignal      => LEDDCLK_ipd,
        RefSignalName  => "LEDDCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_LEDDDAT4_LEDDCLK_posedge_posedge,
        SetupLow       => tsetup_LEDDDAT4_LEDDCLK_negedge_posedge,
        HoldLow        => thold_LEDDDAT4_LEDDCLK_posedge_posedge,
        HoldHigh       => thold_LEDDDAT4_LEDDCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_LEDD_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
		
		
		   VitalSetupHoldCheck (
        Violation      => Tviol_LEDDDAT5_LEDDCLK_posedge,
        TimingData     => Tmkr_LEDDDAT5_LEDDCLK_posedge,
        TestSignal     => LEDDDAT5_ipd,
        TestSignalName => "LEDDDAT5",
        TestDelay      => 0 ns,
        RefSignal      => LEDDCLK_ipd,
        RefSignalName  => "LEDDCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_LEDDDAT5_LEDDCLK_posedge_posedge,
        SetupLow       => tsetup_LEDDDAT5_LEDDCLK_negedge_posedge,
        HoldLow        => thold_LEDDDAT5_LEDDCLK_posedge_posedge,
        HoldHigh       => thold_LEDDDAT5_LEDDCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_LEDD_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
		
		
		   VitalSetupHoldCheck (
        Violation      => Tviol_LEDDDAT6_LEDDCLK_posedge,
        TimingData     => Tmkr_LEDDDAT6_LEDDCLK_posedge,
        TestSignal     => LEDDDAT6_ipd,
        TestSignalName => "LEDDDAT6",
        TestDelay      => 0 ns,
        RefSignal      => LEDDCLK_ipd,
        RefSignalName  => "LEDDCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_LEDDDAT6_LEDDCLK_posedge_posedge,
        SetupLow       => tsetup_LEDDDAT6_LEDDCLK_negedge_posedge,
        HoldLow        => thold_LEDDDAT6_LEDDCLK_posedge_posedge,
        HoldHigh       => thold_LEDDDAT6_LEDDCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_LEDD_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
		
		
		   VitalSetupHoldCheck (
        Violation      => Tviol_LEDDDAT7_LEDDCLK_posedge,
        TimingData     => Tmkr_LEDDDAT7_LEDDCLK_posedge,
        TestSignal     => LEDDDAT7_ipd,
        TestSignalName => "LEDDDAT7",
        TestDelay      => 0 ns,
        RefSignal      => LEDDCLK_ipd,
        RefSignalName  => "LEDDCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_LEDDDAT7_LEDDCLK_posedge_posedge,
        SetupLow       => tsetup_LEDDDAT7_LEDDCLK_negedge_posedge,
        HoldLow        => thold_LEDDDAT7_LEDDCLK_posedge_posedge,
        HoldHigh       => thold_LEDDDAT7_LEDDCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_LEDD_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
end if; 		
----------------------
  --  Path Delay Section
  ----------------------
		
		    VitalPathDelay01 (
      OutSignal     => LEDDON,
      GlitchData    => LEDDON_GlitchData,
      OutSignalName => "LEDDON",
      OutTemp       => LEDDON_zd,
      Paths         => (0 => (LEDDCLK_ipd'last_event, tpd_LEDDCLK_LEDDON_posedge, true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);	
	    VitalPathDelay01 (
      OutSignal     => PWMOUT0,
      GlitchData    => PWMOUT0_GlitchData,
      OutSignalName => "PWMOUT0",
      OutTemp       => PWMOUT0_zd,
      Paths         => (0 => (LEDDCLK_ipd'last_event, tpd_LEDDCLK_PWMOUT0_posedge, true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);
	  
	     VitalPathDelay01 (
      OutSignal     => PWMOUT1,
      GlitchData    => PWMOUT1_GlitchData,
      OutSignalName => "PWMOUT1",
      OutTemp       => PWMOUT1_zd,
      Paths         => (0 => (LEDDCLK_ipd'last_event, tpd_LEDDCLK_PWMOUT1_posedge, true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);
	     VitalPathDelay01 (
      OutSignal     => PWMOUT2,
      GlitchData    => PWMOUT2_GlitchData,
      OutSignalName => "PWMOUT2",
      OutTemp       => PWMOUT2_zd,
      Paths         => (0 => (LEDDCLK_ipd'last_event, tpd_LEDDCLK_PWMOUT2_posedge, true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning); 
	
end process VITALBehavior;
end 	SB_LEDD_IP_V; 

--------------------------------------------------------------
---     	SB_RGB_DRV 		-------
------------------------------------------------

library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;
entity  SB_RGB_DRV  is 
	generic(
		TimingChecksOn : boolean := true;
        Xon            : boolean := false;
        MsgOn          : boolean := false;
		tipd_RGBLEDEN: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_RGB0PWM: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_RGB1PWM: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_RGB2PWM: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_RGBPU: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tpd_RGB0PWM_RGB0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
		tpd_RGB1PWM_RGB1: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tpd_RGB2PWM_RGB2 : VitalDelayType01 := (0.000 ns, 0.000 ns);	
		RGB0_CURRENT: string:="0b000000"; 
		RGB1_CURRENT: string:="0b000000";
		RGB2_CURRENT: string:="0b000000");   
port(
	RGB0: out std_logic;  
	RGB1: out std_logic;
	RGB2: out std_logic;
	RGBLEDEN  :in std_logic;
	RGB0PWM  :in std_logic;
	RGB1PWM:in std_logic;
	RGB2PWM :in std_logic;
    RGBPU : in std_logic
    );
		attribute VITAL_LEVEL0 of			    
    SB_RGB_DRV  : entity is true;
end SB_RGB_DRV ;


architecture SB_RGB_DRV_V of SB_RGB_DRV is
attribute VITAL_LEVEL0 of
    SB_RGB_DRV_V : architecture is true; 
	signal RGBPU_ipd: std_ulogic := 'X';
	signal RGB0PWM_ipd: std_ulogic := 'X';
	signal RGB1PWM_ipd: std_ulogic := 'X';
	signal RGB2PWM_ipd: std_ulogic := 'X';
	signal RGBLEDEN_ipd: std_ulogic := 'X';
	signal RGB0_sig: std_ulogic := 'X';
	signal RGB1_sig: std_ulogic := 'X';
	signal RGB2_sig: std_ulogic := 'X';

component SB_RGB_DRV_CORE 
	GENERIC (RGB0_CURRENT: string:="0b000000"; RGB1_CURRENT: string:="0b000000";RGB2_CURRENT: string:="0b000000");
	port (RGB0: out std_logic;  
	RGB1: out std_logic;
	RGB2: out std_logic;
	RGBLED_EN  :in std_logic;
	RGB0_PWM  :in std_logic;
	RGB1_PWM:in std_logic;
	RGB2_PWM :in std_logic;
    RGB_PU : in std_logic);
end component; 
begin
 WireDelay : block
  begin
    VitalWireDelay (RGBLEDEN_ipd,RGBLEDEN , tipd_RGBLEDEN);
	VitalWireDelay (RGB0PWM_ipd, RGB0PWM, tipd_RGB0PWM);
	VitalWireDelay (RGB1PWM_ipd, RGB0PWM, tipd_RGB1PWM);
	VitalWireDelay (RGB2PWM_ipd, RGB0PWM, tipd_RGB2PWM);
	VitalWireDelay (RGBPU_ipd, RGBPU, tipd_RGBPU);

  end block;
	
LS: SB_RGB_DRV_CORE 
GENERIC MAP (RGB0_CURRENT=>RGB0_CURRENT, RGB1_CURRENT=>RGB1_CURRENT,RGB2_CURRENT=>RGB2_CURRENT)
port map( RGB0=>RGB0_sig,  
	RGB1=>RGB1_sig,
	RGB2=>RGB2_sig ,
	RGBLED_EN=>RGBLEDEN_ipd, 
	RGB0_PWM=>RGB0PWM_ipd, 
	RGB1_PWM=>RGB1PWM_ipd,
	RGB2_PWM=>RGB2PWM_ipd, 
    RGB_PU=>RGBPU_ipd);
VITALPathDelay :process (RGBLEDEN_ipd,RGB0PWM_ipd,RGB1PWM_ipd,RGB2PWM_ipd,RGBPU_ipd,RGB0_sig,RGB1_sig,RGB2_sig)
	variable RGB0_GlitchData : VitalGlitchDataType;
	variable RGB1_GlitchData : VitalGlitchDataType;
	variable RGB2_GlitchData : VitalGlitchDataType;		 
	variable RGB0_zd :std_ulogic:='X'; 
	variable RGB1_zd :std_ulogic:='X';
	variable RGB2_zd :std_ulogic:='X';

		
begin			
	RGB0_zd:=RGB0_sig; 
	RGB1_zd:=RGB1_sig;
	RGB2_zd:=RGB2_sig;
	
VitalPathDelay01 (
      OutSignal                 => RGB0,
      GlitchData                => RGB0_GlitchData,
      OutSignalName             => "RGB0",
      OutTemp                   => RGB0_zd,
      Paths                     => ( 0 =>(RGB0PWM_ipd'last_event, tpd_RGB0PWM_RGB0, true)),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
VitalPathDelay01 (
      OutSignal                 => RGB1,
      GlitchData                => RGB1_GlitchData,
      OutSignalName             => "RGB1",
      OutTemp                   => RGB1_zd,
      Paths                     => (0 =>(RGB1PWM_ipd'last_event, tpd_RGB1PWM_RGB1, true)),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
VitalPathDelay01 (
      OutSignal                 => RGB2,
      GlitchData                => RGB2_GlitchData,
      OutSignalName             => "RGB2",
      OutTemp                   => RGB2_zd,
      Paths                     => (0 =>(RGB2PWM_ipd'last_event, tpd_RGB2PWM_RGB2, true)),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
end process;		 

end 	SB_RGB_DRV_V; 

-------------------------------------------------
---     	SB_LED_DRV_CUR 		-------
------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;
entity SB_LED_DRV_CUR is
	generic( 
		TimingChecksOn : boolean := true;
        Xon            : boolean := false;
        MsgOn          : boolean := false;
		tipd_EN: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tpd_EN_LEDPU : VitalDelayType01 := (0.000 ns, 0.000 ns));
    Port ( EN : in  STD_LOGIC;
           LEDPU : out  STD_LOGIC);
	attribute VITAL_LEVEL0 of			    
    SB_LED_DRV_CUR  : entity is true;
end SB_LED_DRV_CUR;

architecture Behavioral of SB_LED_DRV_CUR is
attribute VITAL_LEVEL0 of
    Behavioral : architecture is true;
	signal EN_ipd: std_ulogic := 'X';
	signal LEDPU_sig: std_ulogic := 'X';
begin
WireDelay : block
  begin
    VitalWireDelay (EN_ipd, EN, tipd_EN);
  end block; 
  process (EN_ipd) 
  begin
  if (EN_ipd = '1') then
	  LEDPU_sig <= '0';
  else
	  LEDPU_sig <= '1';
  end if;	   
  end process;
	--LEDPU_zd <= '0' when (EN_ipd = '1') else '1';
	
VITALPathDelay :process (EN_ipd,LEDPU_sig)
variable LEDPU_GlitchData : VitalGlitchDataType; 
variable LEDPU_zd: std_ulogic := 'X';
begin								 
	   LEDPU_zd:=LEDPU_sig;
VitalPathDelay01 (
      OutSignal                 => LEDPU,
      GlitchData                => LEDPU_GlitchData,
      OutSignalName             => "LEDPU",
      OutTemp                   => LEDPU_zd,
      Paths                     => (0 =>(EN_ipd'last_event, tpd_EN_LEDPU, true)),
      Mode                      => VitalTransport,
      Xon                       => Xon,
      MsgOn                     => MsgOn,
      MsgSeverity               => warning);
end process;
end Behavioral;




-------------------------------------------------
---     	SB_BARCODE_DRV 		-------
------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
use IEEE.VITAL_Timing.all; 
USE IEEE.numeric_std.ALL;
entity  SB_BARCODE_DRV  is
Generic 
(
    TimingChecksOn  : boolean := true;
    Xon   : boolean := true;					   
    MsgOn : boolean := false;
    tpd_BARCODEPWM_BARCODE : VitalDelayType01 := (0 ns, 0 ns);
    tpd_BARCODEEN_BARCODE : VitalDelayType01 := (0 ns, 0 ns);
  	tipd_BARCODEEN 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 	tipd_BARCODEPWM 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 	tipd_CURREN 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
	BARCODE_CURRENT :string := "0b0000";
	CURRENT_MODE :string := "0b0"
);
port (
        BARCODEEN : in std_logic;
		 BARCODEPWM : in std_logic;
		 CURREN : in std_logic;
        BARCODE : out std_logic
	);	 
attribute VITAL_LEVEL0 of
    SB_BARCODE_DRV  : entity is true;
end SB_BARCODE_DRV;

architecture SB_BARCODE_DRV_CORE_V of SB_BARCODE_DRV is
  attribute VITAL_LEVEL0 of
    SB_BARCODE_DRV_CORE_V: architecture is true;

       signal  BARCODEEN_ipd	: std_ulogic :='X' ;
       signal  BARCODEPWM_ipd	: std_ulogic :='X' ;
       signal  CURREN_ipd	: std_ulogic :='X' ;
      signal BARCODE_sig: std_ulogic     := 'X';
	component SB_BARCODE_DRV_CORE
     generic (
		   BARCODE_CURRENT :string := "0b0000";
		    CURRENT_MODE :string := "0b0"
	);
		port ( BARCODEEN : in std_logic;
		 BARCODEPWM : in std_logic;
		 CURREN : in std_logic;
       	 BARCODE : out std_logic
	                	);
	end component;

    begin
    WireDelay:block
    begin
      VitalWireDelay (BARCODEEN_ipd, BARCODEEN, tipd_BARCODEEN);
       VitalWireDelay (BARCODEPWM_ipd, BARCODEPWM, tipd_BARCODEPWM);
       VitalWireDelay (CURREN_ipd, CURREN, tipd_CURREN);

    end block;
		INST: SB_BARCODE_DRV_CORE
		generic map (
			BARCODE_CURRENT =>  BARCODE_CURRENT ,
		    CURRENT_MODE =>  CURRENT_MODE
		)
		port map (
		 BARCODEEN =>  BARCODEEN_ipd   ,
		  BARCODEPWM =>  BARCODEPWM_ipd   ,
		  CURREN =>  CURREN_ipd   ,
       	 BARCODE =>  BARCODE_sig   
		);
VITALPathDelay   : process (  BARCODEEN_ipd, BARCODEPWM_ipd, CURREN_ipd, BARCODE_sig)
variable BARCODE_GlitchData : VitalGlitchDataType;
 variable BARCODE_zd: std_logic :='X';
begin
BARCODE_zd := BARCODE_sig;

     VitalPathDelay01 (
	      OutSignal     => BARCODE,
	      GlitchData    => BARCODE_GlitchData,
	      OutSignalName => "BARCODE",
	      OutTemp       => BARCODE_zd,
	      Paths         => (0 => (BARCODEPWM_ipd'last_event, tpd_BARCODEPWM_BARCODE, true),
							1 => (BARCODEEN_ipd'last_event, tpd_BARCODEEN_BARCODE, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
 end process VITALPathDelay;
end  SB_BARCODE_DRV_CORE_V;		

	


-------------------------------------------------
---     	SB_IR400_DRV 		-------
------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
use IEEE.VITAL_Timing.all; 
USE IEEE.numeric_std.ALL;
entity  SB_IR400_DRV  is
Generic 
(
    TimingChecksOn  : boolean := true;
    Xon   : boolean := true;					   
    MsgOn : boolean := false;
        tpd_IRLEDEN_IRLED : VitalDelayType01 := (0 ns, 0 ns);
       tpd_IRPWM_IRLED : VitalDelayType01 := (0 ns, 0 ns);
  		tipd_CURREN 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_IRLEDEN 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_IRPWM 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
	   CURRENT_MODE :string := "0b0";
		    IR400_CURRENT :string := "0b00000000"
);
port (
        CURREN : in std_logic;
		 IRLEDEN : in std_logic;
		 IRPWM : in std_logic;
        IRLED : out std_logic
	);	 
attribute VITAL_LEVEL0 of
    SB_IR400_DRV  : entity is true;
end SB_IR400_DRV;

architecture SB_IR400_DRV_CORE_V of SB_IR400_DRV is
  attribute VITAL_LEVEL0 of
    SB_IR400_DRV_CORE_V: architecture is true;

          signal  CURREN_ipd	: std_ulogic :='X' ;
       signal  IRLEDEN_ipd	: std_ulogic :='X' ;
       signal  IRPWM_ipd	: std_ulogic :='X' ;

      signal IRLED_sig: std_ulogic     := 'X';
	component SB_IR400_DRV_CORE
     generic (
		   CURRENT_MODE :string := "0b0";
		    IR400_CURRENT :string := "0b00000000"
	);
		port ( CURREN : in std_logic;
		 IRLEDEN : in std_logic;
		 IRPWM : in std_logic;
       			 IRLED : out std_logic
	                	);
	end component;

    begin
    WireDelay:block
    begin
      VitalWireDelay (CURREN_ipd, CURREN, tipd_CURREN);
       VitalWireDelay (IRLEDEN_ipd, IRLEDEN, tipd_IRLEDEN);
       VitalWireDelay (IRPWM_ipd, IRPWM, tipd_IRPWM);

    end block;
		INST: SB_IR400_DRV_CORE
		generic map (
			  CURRENT_MODE =>  CURRENT_MODE ,
		    IR400_CURRENT =>  IR400_CURRENT
		)
		port map (
		 CURREN =>  CURREN_ipd   ,
		  IRLEDEN =>  IRLEDEN_ipd   ,
		  IRPWM =>  IRPWM_ipd   ,
       	 	 IRLED =>  IRLED_sig   
		);
VITALPathDelay   : process (  CURREN_ipd, IRLEDEN_ipd, IRPWM_ipd, IRLED_sig)
variable IRLED_GlitchData : VitalGlitchDataType;
 variable IRLED_zd: std_logic :='X';
begin
IRLED_zd := IRLED_sig;

     VitalPathDelay01 (
	      OutSignal     => IRLED,
	      GlitchData    => IRLED_GlitchData,
	      OutSignalName => "IRLED",
	      OutTemp       => IRLED_zd,
	      Paths         => (0 => (IRLEDEN_ipd'last_event, tpd_IRLEDEN_IRLED, true),
 1 => (IRPWM_ipd'last_event, tpd_IRPWM_IRLED, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
 end process VITALPathDelay;
end  SB_IR400_DRV_CORE_V;		

	



-------------------------------------------------
---     	SB_IR500_DRV 		-------
------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
use IEEE.VITAL_Timing.all; 
USE IEEE.numeric_std.ALL;
entity  SB_IR500_DRV  is
Generic 
(
    TimingChecksOn  : boolean := true;
    Xon   : boolean := true;					   
    MsgOn : boolean := false;
    tpd_IRPWM_IRLED1 : VitalDelayType01 := (0 ns, 0 ns);
    tpd_IRLEDEN_IRLED1 : VitalDelayType01 := (0 ns, 0 ns);
    tpd_IRPWM_IRLED2 : VitalDelayType01 := (0 ns, 0 ns);
    tpd_IRLEDEN_IRLED2 : VitalDelayType01 := (0 ns, 0 ns);
  	tipd_CURREN 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 	tipd_IRLEDEN 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 	tipd_IRPWM 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
	CURRENT_MODE :string := "0b0";
	IR500_CURRENT :string := "0b000000000000"
);
port (
        CURREN : in std_logic;
		IRLEDEN : in std_logic;
		IRPWM : in std_logic;
        IRLED1 : out std_logic;
		IRLED2 : out std_logic
	);	 
attribute VITAL_LEVEL0 of
    SB_IR500_DRV  : entity is true;
end SB_IR500_DRV;

architecture SB_IR500_DRV_CORE_V of SB_IR500_DRV is
  attribute VITAL_LEVEL0 of
    SB_IR500_DRV_CORE_V: architecture is true;

       signal  CURREN_ipd	: std_ulogic :='X' ;
       signal  IRLEDEN_ipd	: std_ulogic :='X' ;
       signal  IRPWM_ipd	: std_ulogic :='X' ;

      signal IRLED1_sig: std_ulogic     := 'X';
      signal IRLED2_sig: std_ulogic     := 'X';
	component SB_IR500_DRV_CORE
     generic (
		   CURRENT_MODE :string := "0b0";
		    IR500_CURRENT :string := "0b000000000000"
	);
		port ( CURREN : in std_logic;
		 IRLEDEN : in std_logic;
		 IRPWM : in std_logic;
       	 IRLED1 : out std_logic;
		 IRLED2 : out std_logic
	                	);
	end component;

    begin
    WireDelay:block
    begin
      VitalWireDelay (CURREN_ipd, CURREN, tipd_CURREN);
       VitalWireDelay (IRLEDEN_ipd, IRLEDEN, tipd_IRLEDEN);
       VitalWireDelay (IRPWM_ipd, IRPWM, tipd_IRPWM);

    end block;
		INST: SB_IR500_DRV_CORE
		generic map (
			CURRENT_MODE =>  CURRENT_MODE ,
		    IR500_CURRENT =>  IR500_CURRENT
		)
		port map (
		 CURREN =>  CURREN_ipd   ,
		  IRLEDEN =>  IRLEDEN_ipd   ,
		  IRPWM =>  IRPWM_ipd   ,
       	  IRLED1 =>  IRLED1_sig   ,
		  IRLED2 =>  IRLED2_sig   
		);
VITALPathDelay   : process ( IRLED1_sig, CURREN_ipd, IRLEDEN_ipd, IRPWM_ipd, IRLED2_sig)
variable IRLED1_GlitchData : VitalGlitchDataType;
 variable IRLED1_zd: std_logic :='X';
 variable IRLED2_GlitchData : VitalGlitchDataType;
 variable IRLED2_zd: std_logic :='X';
begin
IRLED1_zd := IRLED1_sig;
 IRLED2_zd := IRLED2_sig;

     VitalPathDelay01 (
	      OutSignal     => IRLED2,
	      GlitchData    => IRLED2_GlitchData,
	      OutSignalName => "IRLED2",
	      OutTemp       => IRLED2_zd,
	      Paths         => (0 => (IRPWM_ipd'last_event, tpd_IRPWM_IRLED2, true),
							1 => (IRLEDEN_ipd'last_event, tpd_IRLEDEN_IRLED2, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => IRLED1,
	      GlitchData    => IRLED1_GlitchData,
	      OutSignalName => "IRLED1",
	      OutTemp       => IRLED1_zd,
	      Paths         => (0 => (IRPWM_ipd'last_event, tpd_IRPWM_IRLED1, true),
							1 => (IRLEDEN_ipd'last_event, tpd_IRLEDEN_IRLED1, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
 end process VITALPathDelay;
end  SB_IR500_DRV_CORE_V;		



-------------------------------------------------
---     	SB_RGBA_DRV 		-------
------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
use IEEE.VITAL_Timing.all; 
USE IEEE.numeric_std.ALL;
entity  SB_RGBA_DRV  is
Generic 
(
    TimingChecksOn  : boolean := true;
    Xon   : boolean := true;					   
    MsgOn : boolean := false;
        tpd_RGB0PWM_RGB0 : VitalDelayType01 := (0 ns, 0 ns);
       tpd_RGBLEDEN_RGB0 : VitalDelayType01 := (0 ns, 0 ns);
       tpd_RGB1PWM_RGB1 : VitalDelayType01 := (0 ns, 0 ns);
       tpd_RGBLEDEN_RGB1 : VitalDelayType01 := (0 ns, 0 ns);
       tpd_RGB2PWM_RGB2 : VitalDelayType01 := (0 ns, 0 ns);
       tpd_RGBLEDEN_RGB2 : VitalDelayType01 := (0 ns, 0 ns);
  		tipd_CURREN 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_RGB0PWM 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_RGB1PWM 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_RGB2PWM 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_RGBLEDEN 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
	   CURRENT_MODE :string := "0b0";
		    RGB0_CURRENT :string := "0b000000";
		    RGB1_CURRENT :string := "0b000000";
		    RGB2_CURRENT :string := "0b000000"
);
port (
        CURREN : in std_logic;
		 RGB0PWM : in std_logic;
		 RGB1PWM : in std_logic;
		 RGB2PWM : in std_logic;
		 RGBLEDEN : in std_logic;
        RGB0 : out std_logic;
		 RGB1 : out std_logic;
		 RGB2 : out std_logic
	);	 
attribute VITAL_LEVEL0 of
    SB_RGBA_DRV  : entity is true;
end SB_RGBA_DRV;

architecture SB_RGBA_DRV_CORE_V of SB_RGBA_DRV is
  attribute VITAL_LEVEL0 of
    SB_RGBA_DRV_CORE_V: architecture is true;

          signal  CURREN_ipd	: std_ulogic :='X' ;
       signal  RGB0PWM_ipd	: std_ulogic :='X' ;
       signal  RGB1PWM_ipd	: std_ulogic :='X' ;
       signal  RGB2PWM_ipd	: std_ulogic :='X' ;
       signal  RGBLEDEN_ipd	: std_ulogic :='X' ;

      signal RGB0_sig: std_ulogic     := 'X';
        signal RGB1_sig: std_ulogic     := 'X';
        signal RGB2_sig: std_ulogic     := 'X';
	component SB_RGBA_DRV_CORE
     generic (
		   CURRENT_MODE :string := "0b0";
		    RGB0_CURRENT :string := "0b000000";
		    RGB1_CURRENT :string := "0b000000";
		    RGB2_CURRENT :string := "0b000000"
	);
		port ( CURREN : in std_logic;
		 RGB0PWM : in std_logic;
		 RGB1PWM : in std_logic;
		 RGB2PWM : in std_logic;
		 RGBLEDEN : in std_logic;
       			 RGB0 : out std_logic;
		 RGB1 : out std_logic;
		 RGB2 : out std_logic
	                	);
	end component;

    begin
    WireDelay:block
    begin
      VitalWireDelay (CURREN_ipd, CURREN, tipd_CURREN);
       VitalWireDelay (RGB0PWM_ipd, RGB0PWM, tipd_RGB0PWM);
       VitalWireDelay (RGB1PWM_ipd, RGB1PWM, tipd_RGB1PWM);
       VitalWireDelay (RGB2PWM_ipd, RGB2PWM, tipd_RGB2PWM);
       VitalWireDelay (RGBLEDEN_ipd, RGBLEDEN, tipd_RGBLEDEN);

    end block;
		INST: SB_RGBA_DRV_CORE
		generic map (
			  CURRENT_MODE =>  CURRENT_MODE ,
		   RGB0_CURRENT =>  RGB0_CURRENT ,
		   RGB1_CURRENT =>  RGB1_CURRENT ,
		    RGB2_CURRENT =>  RGB2_CURRENT
		)
		port map (
		 CURREN =>  CURREN_ipd   ,
		  RGB0PWM =>  RGB0PWM_ipd   ,
		  RGB1PWM =>  RGB1PWM_ipd   ,
		  RGB2PWM =>  RGB2PWM_ipd   ,
		  RGBLEDEN =>  RGBLEDEN_ipd   ,
       	 	 RGB0 =>  RGB0_sig   ,
		  RGB1 =>  RGB1_sig   ,
		  RGB2 =>  RGB2_sig   
		);
VITALPathDelay   : process ( RGB0_sig, RGB1_sig, CURREN_ipd, RGB0PWM_ipd, RGB1PWM_ipd, RGB2PWM_ipd, RGBLEDEN_ipd, RGB2_sig)
variable RGB0_GlitchData : VitalGlitchDataType;
 variable RGB0_zd: std_logic :='X';
 variable RGB1_GlitchData : VitalGlitchDataType;
 variable RGB1_zd: std_logic :='X';
 variable RGB2_GlitchData : VitalGlitchDataType;
 variable RGB2_zd: std_logic :='X';
begin
RGB0_zd := RGB0_sig;
 RGB1_zd := RGB1_sig;
 RGB2_zd := RGB2_sig;

     VitalPathDelay01 (
	      OutSignal     => RGB0,
	      GlitchData    => RGB0_GlitchData,
	      OutSignalName => "RGB0",
	      OutTemp       => RGB0_zd,
	      Paths         => (0 => (RGB0PWM_ipd'last_event, tpd_RGB0PWM_RGB0, true),
 1 => (RGBLEDEN_ipd'last_event, tpd_RGBLEDEN_RGB0, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => RGB1,
	      GlitchData    => RGB1_GlitchData,
	      OutSignalName => "RGB1",
	      OutTemp       => RGB1_zd,
	      Paths         => (0 => (RGB1PWM_ipd'last_event, tpd_RGB1PWM_RGB1, true),
 1 => (RGBLEDEN_ipd'last_event, tpd_RGBLEDEN_RGB1, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => RGB2,
	      GlitchData    => RGB2_GlitchData,
	      OutSignalName => "RGB2",
	      OutTemp       => RGB2_zd,
	      Paths         => (0 => (RGB2PWM_ipd'last_event, tpd_RGB2PWM_RGB2, true),
 1 => (RGBLEDEN_ipd'last_event, tpd_RGBLEDEN_RGB2, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
 end process VITALPathDelay;
end  SB_RGBA_DRV_CORE_V;		




-------------------------------------------------
---     	SB_I2C_FIFO 		-------
------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
use IEEE.VITAL_Timing.all; 
USE IEEE.numeric_std.ALL;
entity  SB_I2C_FIFO  is
Generic 
(
    TimingChecksOn  : boolean := true;
    Xon   : boolean := true;					   
    MsgOn : boolean := false;
	
		tsetup_SDAI_SCLO_negedge_posedge : VitalDelayType := 0 ns;
 		tsetup_SDAI_SCLO_posedge_posedge : VitalDelayType:= 0 ns;
 		thold_SDAI_SCLO_negedge_posedge : VitalDelayType := 0 ns;
 		thold_SDAI_SCLO_posedge_posedge : VitalDelayType:= 0 ns;
		tsetup_SDAI_SCLI_negedge_posedge : VitalDelayType := 0 ns;
 		tsetup_SDAI_SCLI_posedge_posedge : VitalDelayType:= 0 ns;
 		thold_SDAI_SCLI_negedge_posedge : VitalDelayType := 0 ns;
 		thold_SDAI_SCLI_posedge_posedge : VitalDelayType:= 0 ns;
  		tsetup_CSI_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		tsetup_CSI_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		thold_CSI_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		thold_CSI_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		tsetup_STBI_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		tsetup_STBI_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		thold_STBI_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		thold_STBI_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		tsetup_WEI_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		tsetup_WEI_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		thold_WEI_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		thold_WEI_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		tsetup_FIFORST_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		tsetup_FIFORST_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		thold_FIFORST_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		thold_FIFORST_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		tsetup_SDAI_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		tsetup_SDAI_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		thold_SDAI_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		thold_SDAI_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		tsetup_ADRI3_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		tsetup_ADRI3_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		thold_ADRI3_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		thold_ADRI3_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		tsetup_ADRI2_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		tsetup_ADRI2_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		thold_ADRI2_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		thold_ADRI2_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		tsetup_ADRI1_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		tsetup_ADRI1_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		thold_ADRI1_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		thold_ADRI1_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		tsetup_ADRI0_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		tsetup_ADRI0_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		thold_ADRI0_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		thold_ADRI0_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		tsetup_DATI0_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		tsetup_DATI0_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		thold_DATI0_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		thold_DATI0_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		tsetup_DATI1_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		tsetup_DATI1_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		thold_DATI1_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		thold_DATI1_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		tsetup_DATI2_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		tsetup_DATI2_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		thold_DATI2_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		thold_DATI2_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		tsetup_DATI3_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		tsetup_DATI3_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		thold_DATI3_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		thold_DATI3_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		tsetup_DATI4_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		tsetup_DATI4_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		thold_DATI4_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		thold_DATI4_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		tsetup_DATI5_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		tsetup_DATI5_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		thold_DATI5_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		thold_DATI5_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		tsetup_DATI6_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		tsetup_DATI6_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		thold_DATI6_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		thold_DATI6_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		tsetup_DATI7_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		tsetup_DATI7_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		thold_DATI7_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		thold_DATI7_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		tsetup_DATI8_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		tsetup_DATI8_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		thold_DATI8_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		thold_DATI8_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		tsetup_DATI9_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		tsetup_DATI9_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		thold_DATI9_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		thold_DATI9_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		tsetup_SCLO_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		tsetup_SCLO_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		thold_SCLO_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		thold_SCLO_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		tsetup_SCLI_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		tsetup_SCLI_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
 		thold_SCLI_CLKI_negedge_posedge : VitalDelayType := 0 ns;
 		thold_SCLI_CLKI_posedge_posedge : VitalDelayType:= 0 ns;

  		tpw_CLKI_posedge : VitalDelayType := 0 ns;
 		tpw_CLKI_negedge : VitalDelayType := 0 ns;

  		tpd_CLKI_SCLO : VitalDelayType01 := (0 ns, 0 ns);
 		 tpd_CLKI_SCLO_posedge : VitalDelayType01 := (0 ns, 0 ns);
 		tpd_CLKI_ACKO : VitalDelayType01 := (0 ns, 0 ns);
 		 tpd_CLKI_ACKO_posedge : VitalDelayType01 := (0 ns, 0 ns);
 		tpd_CLKI_DATO0 : VitalDelayType01 := (0 ns, 0 ns);
 		 tpd_CLKI_DATO0_posedge : VitalDelayType01 := (0 ns, 0 ns);
 		tpd_CLKI_DATO1 : VitalDelayType01 := (0 ns, 0 ns);
 		 tpd_CLKI_DATO1_posedge : VitalDelayType01 := (0 ns, 0 ns);
 		tpd_CLKI_DATO2 : VitalDelayType01 := (0 ns, 0 ns);
 		 tpd_CLKI_DATO2_posedge : VitalDelayType01 := (0 ns, 0 ns);
 		tpd_CLKI_DATO3 : VitalDelayType01 := (0 ns, 0 ns);
 		 tpd_CLKI_DATO3_posedge : VitalDelayType01 := (0 ns, 0 ns);
 		tpd_CLKI_DATO4 : VitalDelayType01 := (0 ns, 0 ns);
 		 tpd_CLKI_DATO4_posedge : VitalDelayType01 := (0 ns, 0 ns);
 		tpd_CLKI_DATO5 : VitalDelayType01 := (0 ns, 0 ns);
 		 tpd_CLKI_DATO5_posedge : VitalDelayType01 := (0 ns, 0 ns);
 		tpd_CLKI_DATO6 : VitalDelayType01 := (0 ns, 0 ns);
 		 tpd_CLKI_DATO6_posedge : VitalDelayType01 := (0 ns, 0 ns);
 		tpd_CLKI_DATO7 : VitalDelayType01 := (0 ns, 0 ns);
 		 tpd_CLKI_DATO7_posedge : VitalDelayType01 := (0 ns, 0 ns);
 		tpd_CLKI_DATO8 : VitalDelayType01 := (0 ns, 0 ns);
 		 tpd_CLKI_DATO8_posedge : VitalDelayType01 := (0 ns, 0 ns);
 		tpd_CLKI_DATO9 : VitalDelayType01 := (0 ns, 0 ns);
 		 tpd_CLKI_DATO9_posedge : VitalDelayType01 := (0 ns, 0 ns);
 		tpd_CLKI_I2CIRQ : VitalDelayType01 := (0 ns, 0 ns);
 		 tpd_CLKI_I2CIRQ_posedge : VitalDelayType01 := (0 ns, 0 ns);
 		tpd_CLKI_I2CWKUP : VitalDelayType01 := (0 ns, 0 ns);
 		 tpd_CLKI_I2CWKUP_posedge : VitalDelayType01 := (0 ns, 0 ns);
 		tpd_CLKI_SCLOE : VitalDelayType01 := (0 ns, 0 ns);
 		 tpd_CLKI_SCLOE_posedge : VitalDelayType01 := (0 ns, 0 ns);
 		tpd_CLKI_SDAO : VitalDelayType01 := (0 ns, 0 ns);
 		 tpd_CLKI_SDAO_posedge : VitalDelayType01 := (0 ns, 0 ns);
 		tpd_SCLO_SDAO_posedge : VitalDelayType01 := (0 ns, 0 ns);
        	tpd_SCLO_SDAO_negedge : VitalDelayType01 := (0 ns, 0 ns);
			tpd_SCLI_SDAO_posedge : VitalDelayType01 := (0 ns, 0 ns);
        	tpd_SCLI_SDAO_negedge : VitalDelayType01 := (0 ns, 0 ns);
 		 --tpd_CLKI_SDAO_posedge : VitalDelayType01 := (0 ns, 0 ns);
 		tpd_CLKI_SDAOE : VitalDelayType01 := (0 ns, 0 ns);
 		 tpd_CLKI_SDAOE_posedge : VitalDelayType01 := (0 ns, 0 ns);
 		tpd_SCLO_SDAOE_posedge : VitalDelayType01 := (0 ns, 0 ns);
        	tpd_SCLO_SDAOE_negedge : VitalDelayType01 := (0 ns, 0 ns);
			tpd_SCLI_SDAOE_posedge : VitalDelayType01 := (0 ns, 0 ns);
        	tpd_SCLI_SDAOE_negedge : VitalDelayType01 := (0 ns, 0 ns);
 		 --tpd_CLKI_SDAOE_posedge : VitalDelayType01 := (0 ns, 0 ns);
 		tpd_CLKI_SRWO : VitalDelayType01 := (0 ns, 0 ns);
 		 tpd_CLKI_SRWO_posedge : VitalDelayType01 := (0 ns, 0 ns);
 		 
         tpd_CLKI_TXFIFOEMPTY_posedge : VitalDelayType01 := (0 ns, 0 ns);
         tpd_CLKI_TXFIFOAEMPTY_posedge : VitalDelayType01 := (0 ns, 0 ns);
         tpd_CLKI_TXFIFOFULL_posedge : VitalDelayType01 := (0 ns, 0 ns);

         tpd_CLKI_RXFIFOEMPTY_posedge : VitalDelayType01 := (0 ns, 0 ns);
         tpd_CLKI_RXFIFOAFULL_posedge : VitalDelayType01 := (0 ns, 0 ns);
         tpd_CLKI_RXFIFOFULL_posedge : VitalDelayType01 := (0 ns, 0 ns);

         tpd_CLKI_TXFIFOEMPTY_negedge : VitalDelayType01 := (0 ns, 0 ns);
         tpd_CLKI_TXFIFOAEMPTY_negedge : VitalDelayType01 := (0 ns, 0 ns);
         tpd_CLKI_TXFIFOFULL_negedge : VitalDelayType01 := (0 ns, 0 ns);

         tpd_CLKI_RXFIFOEMPTY_negedge : VitalDelayType01 := (0 ns, 0 ns);
         tpd_CLKI_RXFIFOAFULL_negedge : VitalDelayType01 := (0 ns, 0 ns);
         tpd_CLKI_RXFIFOFULL_negedge : VitalDelayType01 := (0 ns, 0 ns);

  		I2C_SLAVE_ADDR :string := "0b1111100001";

  		tipd_ADRI0 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_ADRI1 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_ADRI2 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_ADRI3 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_CLKI 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_CSI 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_DATI0 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_DATI1 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_DATI2 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_DATI3 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_DATI4 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_DATI5 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_DATI6 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_DATI7 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_DATI8 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_DATI9 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_FIFORST 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_SCLI 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_SDAI 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_STBI 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_SCLO 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_WEI 	: VitalDelayType01 := (0.000 ns, 0.000 ns)
);
port (
        ADRI0 : in std_logic;
		 ADRI1 : in std_logic;
		 ADRI2 : in std_logic;
		 ADRI3 : in std_logic;
		 CLKI : in std_logic;
		 CSI : in std_logic;
		 DATI0 : in std_logic :='L';
		 DATI1 : in std_logic :='L';
		 DATI2 : in std_logic :='L';
		 DATI3 : in std_logic :='L';
		 DATI4 : in std_logic :='L';
		 DATI5 : in std_logic :='L';
		 DATI6 : in std_logic :='L';
		 DATI7 : in std_logic :='L';
		 DATI8 : in std_logic :='L';
		 DATI9 : in std_logic :='L';
		 FIFORST : in std_logic;
		 SCLI : in std_logic;
		 SDAI : in std_logic;
		 STBI : in std_logic;
		 WEI : in std_logic;
		SCLO : out std_logic;
        ACKO : out std_logic;
		 DATO0 : out std_logic;
		 DATO1 : out std_logic;
		 DATO2 : out std_logic;
		 DATO3 : out std_logic;
		 DATO4 : out std_logic;
		 DATO5 : out std_logic;
		 DATO6 : out std_logic;
		 DATO7 : out std_logic;
		 DATO8 : out std_logic;
		 DATO9 : out std_logic;
		 I2CIRQ : out std_logic;
		 I2CWKUP : out std_logic;
		 MRDCMPL : out std_logic;
		 RXFIFOAFULL : out std_logic;
		 RXFIFOEMPTY : out std_logic;
		 RXFIFOFULL : out std_logic;
		 SCLOE : out std_logic;
		 SDAO : out std_logic;
		 SDAOE : out std_logic;
		 SRWO : out std_logic;
		 TXFIFOAEMPTY : out std_logic;
		 TXFIFOEMPTY : out std_logic;
		 TXFIFOFULL : out std_logic
	);	 
attribute VITAL_LEVEL0 of
    SB_I2C_FIFO  : entity is true;
end SB_I2C_FIFO;

architecture SB_I2C_FIFO_V of SB_I2C_FIFO is
  attribute VITAL_LEVEL0 of
    SB_I2C_FIFO_V: architecture is true;

    		signal  ADRI0_ipd	: std_ulogic :='X' ;
 		signal  ADRI1_ipd	: std_ulogic :='X' ;
 		signal  ADRI2_ipd	: std_ulogic :='X' ;
 		signal  ADRI3_ipd	: std_ulogic :='X' ;
 		signal  CLKI_ipd	: std_ulogic :='X' ;
 		signal  CSI_ipd	: std_ulogic :='X' ;
 		signal  DATI0_ipd	: std_ulogic :='X' ;
 		signal  DATI1_ipd	: std_ulogic :='X' ;
 		signal  DATI2_ipd	: std_ulogic :='X' ;
 		signal  DATI3_ipd	: std_ulogic :='X' ;
 		signal  DATI4_ipd	: std_ulogic :='X' ;
 		signal  DATI5_ipd	: std_ulogic :='X' ;
 		signal  DATI6_ipd	: std_ulogic :='X' ;
 		signal  DATI7_ipd	: std_ulogic :='X' ;
 		signal  DATI8_ipd	: std_ulogic :='X' ;
 		signal  DATI9_ipd	: std_ulogic :='X' ;
 		signal  FIFORST_ipd	: std_ulogic :='X' ;
 		signal  SCLI_ipd	: std_ulogic :='X' ;
 		signal  SDAI_ipd	: std_ulogic :='X' ;
 		signal  STBI_ipd	: std_ulogic :='X' ;
 		signal  WEI_ipd	: std_ulogic :='X' ;
		signal  SCLO_ipd	: std_ulogic :='X' ;
		signal SCLO_sig: std_ulogic     := 'X';
		signal ACKO_sig: std_ulogic     := 'X';
  		signal DATO0_sig: std_ulogic     := 'X';
  		signal DATO1_sig: std_ulogic     := 'X';
  		signal DATO2_sig: std_ulogic     := 'X';
  		signal DATO3_sig: std_ulogic     := 'X';
  		signal DATO4_sig: std_ulogic     := 'X';
  		signal DATO5_sig: std_ulogic     := 'X';
  		signal DATO6_sig: std_ulogic     := 'X';
  		signal DATO7_sig: std_ulogic     := 'X';
  		signal DATO8_sig: std_ulogic     := 'X';
  		signal DATO9_sig: std_ulogic     := 'X';
  		signal I2CIRQ_sig: std_ulogic     := 'X';
  		signal I2CWKUP_sig: std_ulogic     := 'X';
  		signal MRDCMPL_sig: std_ulogic     := 'X';
  		signal RXFIFOAFULL_sig: std_ulogic     := 'X';
  		signal RXFIFOEMPTY_sig: std_ulogic     := 'X';
  		signal RXFIFOFULL_sig: std_ulogic     := 'X';
  		signal SCLOE_sig: std_ulogic     := 'X';
  		signal SDAO_sig: std_ulogic     := 'X';
  		signal SDAOE_sig: std_ulogic     := 'X';
  		signal SRWO_sig: std_ulogic     := 'X';
  		signal TXFIFOAEMPTY_sig: std_ulogic     := 'X';
  		signal TXFIFOEMPTY_sig: std_ulogic     := 'X';
  		signal TXFIFOFULL_sig: std_ulogic     := 'X';
	component SB_I2C_FIFO_CORE
     generic (
				I2C_SLAVE_ADDR :string := "0b1111100001"
	);
		port ( 
		ADRI0 : in std_logic;
		 ADRI1 : in std_logic;
		 ADRI2 : in std_logic;
		 ADRI3 : in std_logic;
		 CLKI : in std_logic;
		 CSI : in std_logic;
		 DATI0 : in std_logic;
		 DATI1 : in std_logic;
		 DATI2 : in std_logic;
		 DATI3 : in std_logic;
		 DATI4 : in std_logic;
		 DATI5 : in std_logic;
		 DATI6 : in std_logic;
		 DATI7 : in std_logic;
		 DATI8 : in std_logic;
		 DATI9 : in std_logic;
		 FIFORST : in std_logic;
		 SCLI : in std_logic;
		 SDAI : in std_logic;
		 STBI : in std_logic;
		 WEI : in std_logic;
		SCLO : out std_logic;
		ACKO : out std_logic;
		 DATO0 : out std_logic;
		 DATO1 : out std_logic;
		 DATO2 : out std_logic;
		 DATO3 : out std_logic;
		 DATO4 : out std_logic;
		 DATO5 : out std_logic;
		 DATO6 : out std_logic;
		 DATO7 : out std_logic;
		 DATO8 : out std_logic;
		 DATO9 : out std_logic;
		 I2CIRQ : out std_logic;
		 I2CWKUP : out std_logic;
		 MRDCMPL : out std_logic;
		 RXFIFOAFULL : out std_logic;
		 RXFIFOEMPTY : out std_logic;
		 RXFIFOFULL : out std_logic;
		 SCLOE : out std_logic;
		 SDAO : out std_logic;
		 SDAOE : out std_logic;
		 SRWO : out std_logic;
		 TXFIFOAEMPTY : out std_logic;
		 TXFIFOEMPTY : out std_logic;
		 TXFIFOFULL : out std_logic
	                	);
	end component;

    begin
    WireDelay:block
    begin
		VitalWireDelay (ADRI0_ipd, ADRI0, tipd_ADRI0);
 		VitalWireDelay (ADRI1_ipd, ADRI1, tipd_ADRI1);
 		VitalWireDelay (ADRI2_ipd, ADRI2, tipd_ADRI2);
 		VitalWireDelay (ADRI3_ipd, ADRI3, tipd_ADRI3);
 		VitalWireDelay (CLKI_ipd, CLKI, tipd_CLKI);
 		VitalWireDelay (CSI_ipd, CSI, tipd_CSI);
 		VitalWireDelay (DATI0_ipd, DATI0, tipd_DATI0);
 		VitalWireDelay (DATI1_ipd, DATI1, tipd_DATI1);
 		VitalWireDelay (DATI2_ipd, DATI2, tipd_DATI2);
 		VitalWireDelay (DATI3_ipd, DATI3, tipd_DATI3);
 		VitalWireDelay (DATI4_ipd, DATI4, tipd_DATI4);
 		VitalWireDelay (DATI5_ipd, DATI5, tipd_DATI5);
 		VitalWireDelay (DATI6_ipd, DATI6, tipd_DATI6);
 		VitalWireDelay (DATI7_ipd, DATI7, tipd_DATI7);
 		VitalWireDelay (DATI8_ipd, DATI8, tipd_DATI8);
 		VitalWireDelay (DATI9_ipd, DATI9, tipd_DATI9);
 		VitalWireDelay (FIFORST_ipd, FIFORST, tipd_FIFORST);
 		VitalWireDelay (SCLI_ipd, SCLI, tipd_SCLI);
 		VitalWireDelay (SDAI_ipd, SDAI, tipd_SDAI);
 		VitalWireDelay (STBI_ipd, STBI, tipd_STBI);
 		VitalWireDelay (WEI_ipd, WEI, tipd_WEI);


    end block;
		INST: SB_I2C_FIFO_CORE
		generic map (
				I2C_SLAVE_ADDR =>  I2C_SLAVE_ADDR
		)
		port map (
		ADRI0 =>  ADRI0_ipd   ,
		 ADRI1 =>  ADRI1_ipd   ,
		 ADRI2 =>  ADRI2_ipd   ,
		 ADRI3 =>  ADRI3_ipd   ,
		 CLKI =>  CLKI_ipd   ,
		 CSI =>  CSI_ipd   ,
		 DATI0 =>  DATI0_ipd   ,
		 DATI1 =>  DATI1_ipd   ,
		 DATI2 =>  DATI2_ipd   ,
		 DATI3 =>  DATI3_ipd   ,
		 DATI4 =>  DATI4_ipd   ,
		 DATI5 =>  DATI5_ipd   ,
		 DATI6 =>  DATI6_ipd   ,
		 DATI7 =>  DATI7_ipd   ,
		 DATI8 =>  DATI8_ipd   ,
		 DATI9 =>  DATI9_ipd   ,
		 FIFORST =>  FIFORST_ipd   ,
		 SCLI =>  SCLI_ipd   ,
		 SDAI =>  SDAI_ipd   ,
		 STBI =>  STBI_ipd   ,
		 WEI =>  WEI_ipd   ,
		 SCLO =>  SCLO_sig   ,
       	 ACKO =>  ACKO_sig   ,
		  DATO0 =>  DATO0_sig   ,
		  DATO1 =>  DATO1_sig   ,
		  DATO2 =>  DATO2_sig   ,
		  DATO3 =>  DATO3_sig   ,
		  DATO4 =>  DATO4_sig   ,
		  DATO5 =>  DATO5_sig   ,
		  DATO6 =>  DATO6_sig   ,
		  DATO7 =>  DATO7_sig   ,
		  DATO8 =>  DATO8_sig   ,
		  DATO9 =>  DATO9_sig   ,
		  I2CIRQ =>  I2CIRQ_sig   ,
		  I2CWKUP =>  I2CWKUP_sig   ,
		  MRDCMPL =>  MRDCMPL_sig   ,
		  RXFIFOAFULL =>  RXFIFOAFULL_sig   ,
		  RXFIFOEMPTY =>  RXFIFOEMPTY_sig   ,
		  RXFIFOFULL =>  RXFIFOFULL_sig   ,
		  SCLOE =>  SCLOE_sig   ,
		  SDAO =>  SDAO_sig   ,
		  SDAOE =>  SDAOE_sig   ,
		  SRWO =>  SRWO_sig   ,
		  TXFIFOAEMPTY =>  TXFIFOAEMPTY_sig   ,
		  TXFIFOEMPTY =>  TXFIFOEMPTY_sig   ,
		  TXFIFOFULL =>  TXFIFOFULL_sig   
		);
VITALBehavior   : process ( SCLO_sig, ACKO_sig, DATO0_sig, DATO1_sig, DATO2_sig, DATO3_sig, DATO4_sig, DATO5_sig, DATO6_sig, DATO7_sig, DATO8_sig, DATO9_sig, I2CIRQ_sig, I2CWKUP_sig, MRDCMPL_sig, RXFIFOAFULL_sig, RXFIFOEMPTY_sig, RXFIFOFULL_sig, SCLOE_sig, SDAO_sig, SDAOE_sig, SRWO_sig, TXFIFOAEMPTY_sig, TXFIFOEMPTY_sig, ADRI0_ipd, ADRI1_ipd, ADRI2_ipd, ADRI3_ipd, CLKI_ipd,SCLO_ipd,SCLI_ipd, CSI_ipd, DATI0_ipd, DATI1_ipd, DATI2_ipd, DATI3_ipd, DATI4_ipd, DATI5_ipd, DATI6_ipd, DATI7_ipd, DATI8_ipd, DATI9_ipd, FIFORST_ipd, SCLI_ipd, SDAI_ipd, STBI_ipd, WEI_ipd,TXFIFOFULL_sig)

		variable      Tviol_CSI_CLKI_posedge : std_logic := '0';
 		variable      Tmkr_CSI_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
 		variable      Tviol_STBI_CLKI_posedge : std_logic := '0';
 		variable      Tmkr_STBI_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
 		variable      Tviol_WEI_CLKI_posedge : std_logic := '0';
 		variable      Tmkr_WEI_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
 		variable      Tviol_FIFORST_CLKI_posedge : std_logic := '0';
 		variable      Tmkr_FIFORST_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
 		variable      Tviol_SDAI_CLKI_posedge : std_logic := '0';
 		variable      Tmkr_SDAI_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
 		variable      Tviol_ADRI3_CLKI_posedge : std_logic := '0';
 		variable      Tmkr_ADRI3_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
 		variable      Tviol_ADRI2_CLKI_posedge : std_logic := '0';
 		variable      Tmkr_ADRI2_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
 		variable      Tviol_ADRI1_CLKI_posedge : std_logic := '0';
 		variable      Tmkr_ADRI1_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
 		variable      Tviol_ADRI0_CLKI_posedge : std_logic := '0';
 		variable      Tmkr_ADRI0_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
 		variable      Tviol_DATI0_CLKI_posedge : std_logic := '0';
 		variable      Tmkr_DATI0_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
 		variable      Tviol_DATI1_CLKI_posedge : std_logic := '0';
 		variable      Tmkr_DATI1_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
 		variable      Tviol_DATI2_CLKI_posedge : std_logic := '0';
 		variable      Tmkr_DATI2_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
 		variable      Tviol_DATI3_CLKI_posedge : std_logic := '0';
 		variable      Tmkr_DATI3_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
 		variable      Tviol_DATI4_CLKI_posedge : std_logic := '0';
 		variable      Tmkr_DATI4_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
 		variable      Tviol_DATI5_CLKI_posedge : std_logic := '0';
 		variable      Tmkr_DATI5_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
 		variable      Tviol_DATI6_CLKI_posedge : std_logic := '0';
 		variable      Tmkr_DATI6_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
 		variable      Tviol_DATI7_CLKI_posedge : std_logic := '0';
 		variable      Tmkr_DATI7_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
 		variable      Tviol_DATI8_CLKI_posedge : std_logic := '0';
 		variable      Tmkr_DATI8_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
 		variable      Tviol_DATI9_CLKI_posedge : std_logic := '0';
 		variable      Tmkr_DATI9_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
 		variable      Tviol_SCLO_CLKI_posedge : std_logic := '0';
 		variable      Tmkr_SCLO_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
 		variable      Tviol_SCLI_CLKI_posedge : std_logic := '0';
 		variable      Tmkr_SCLI_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
		variable      Tviol_SDAI_SCLO_posedge : std_logic := '0';
 		variable      Tmkr_SDAI_SCLO_posedge : VitalTimingDataType :=VitalTimingDataInit ;
		variable      Tviol_SDAI_SCLI_posedge : std_logic := '0';
 		variable      Tmkr_SDAI_SCLI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
variable      Pviol_CLKI : std_logic := '0';
 variable      PInfo_CLKI : VitalPeriodDataType := VitalPeriodDataInit;
begin
if (TimingChecksOn) then
VitalSetupHoldCheck (
        Violation      =>Tviol_SDAI_SCLO_posedge ,
        TimingData     =>Tmkr_SDAI_SCLO_posedge  ,
        TestSignal     => SDAI_ipd,
        TestSignalName => "SDAI",
        TestDelay      => 0 ns,
        RefSignal      => SCLO_ipd,
        RefSignalName  => "SCLO",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_SDAI_SCLO_posedge_posedge ,
        SetupLow       => tsetup_SDAI_SCLO_negedge_posedge,
        HoldLow        => thold_SDAI_SCLO_posedge_posedge,
        HoldHigh       => thold_SDAI_SCLO_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C_FIFO",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
		
VitalSetupHoldCheck (
        Violation      =>Tviol_SDAI_SCLI_posedge ,
        TimingData     =>Tmkr_SDAI_SCLI_posedge  ,
        TestSignal     => SDAI_ipd,
        TestSignalName => "SDAI",
        TestDelay      => 0 ns,
        RefSignal      => SCLI_ipd,
        RefSignalName  => "SCLI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_SDAI_SCLI_posedge_posedge ,
        SetupLow       => tsetup_SDAI_SCLI_negedge_posedge,
        HoldLow        => thold_SDAI_SCLI_posedge_posedge,
        HoldHigh       => thold_SDAI_SCLI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C_FIFO",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	

 VitalSetupHoldCheck (
        Violation      =>Tviol_CSI_CLKI_posedge ,
        TimingData     =>Tmkr_CSI_CLKI_posedge  ,
        TestSignal     => CSI_ipd,
        TestSignalName => "CSI",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_CSI_CLKI_posedge_posedge ,
        SetupLow       => tsetup_CSI_CLKI_negedge_posedge,
        HoldLow        => thold_CSI_CLKI_posedge_posedge,
        HoldHigh       => thold_CSI_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C_FIFO",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_STBI_CLKI_posedge ,
        TimingData     =>Tmkr_STBI_CLKI_posedge  ,
        TestSignal     => STBI_ipd,
        TestSignalName => "STBI",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_STBI_CLKI_posedge_posedge ,
        SetupLow       => tsetup_STBI_CLKI_negedge_posedge,
        HoldLow        => thold_STBI_CLKI_posedge_posedge,
        HoldHigh       => thold_STBI_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C_FIFO",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_WEI_CLKI_posedge ,
        TimingData     =>Tmkr_WEI_CLKI_posedge  ,
        TestSignal     => WEI_ipd,
        TestSignalName => "WEI",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WEI_CLKI_posedge_posedge ,
        SetupLow       => tsetup_WEI_CLKI_negedge_posedge,
        HoldLow        => thold_WEI_CLKI_posedge_posedge,
        HoldHigh       => thold_WEI_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C_FIFO",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_FIFORST_CLKI_posedge ,
        TimingData     =>Tmkr_FIFORST_CLKI_posedge  ,
        TestSignal     => FIFORST_ipd,
        TestSignalName => "FIFORST",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_FIFORST_CLKI_posedge_posedge ,
        SetupLow       => tsetup_FIFORST_CLKI_negedge_posedge,
        HoldLow        => thold_FIFORST_CLKI_posedge_posedge,
        HoldHigh       => thold_FIFORST_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C_FIFO",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_SDAI_CLKI_posedge ,
        TimingData     =>Tmkr_SDAI_CLKI_posedge  ,
        TestSignal     => SDAI_ipd,
        TestSignalName => "SDAI",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_SDAI_CLKI_posedge_posedge ,
        SetupLow       => tsetup_SDAI_CLKI_negedge_posedge,
        HoldLow        => thold_SDAI_CLKI_posedge_posedge,
        HoldHigh       => thold_SDAI_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C_FIFO",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_ADRI3_CLKI_posedge ,
        TimingData     =>Tmkr_ADRI3_CLKI_posedge  ,
        TestSignal     => ADRI3_ipd,
        TestSignalName => "ADRI3",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_ADRI3_CLKI_posedge_posedge ,
        SetupLow       => tsetup_ADRI3_CLKI_negedge_posedge,
        HoldLow        => thold_ADRI3_CLKI_posedge_posedge,
        HoldHigh       => thold_ADRI3_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C_FIFO",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_ADRI2_CLKI_posedge ,
        TimingData     =>Tmkr_ADRI2_CLKI_posedge  ,
        TestSignal     => ADRI2_ipd,
        TestSignalName => "ADRI2",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_ADRI2_CLKI_posedge_posedge ,
        SetupLow       => tsetup_ADRI2_CLKI_negedge_posedge,
        HoldLow        => thold_ADRI2_CLKI_posedge_posedge,
        HoldHigh       => thold_ADRI2_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C_FIFO",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_ADRI1_CLKI_posedge ,
        TimingData     =>Tmkr_ADRI1_CLKI_posedge  ,
        TestSignal     => ADRI1_ipd,
        TestSignalName => "ADRI1",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_ADRI1_CLKI_posedge_posedge ,
        SetupLow       => tsetup_ADRI1_CLKI_negedge_posedge,
        HoldLow        => thold_ADRI1_CLKI_posedge_posedge,
        HoldHigh       => thold_ADRI1_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C_FIFO",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_ADRI0_CLKI_posedge ,
        TimingData     =>Tmkr_ADRI0_CLKI_posedge  ,
        TestSignal     => ADRI0_ipd,
        TestSignalName => "ADRI0",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_ADRI0_CLKI_posedge_posedge ,
        SetupLow       => tsetup_ADRI0_CLKI_negedge_posedge,
        HoldLow        => thold_ADRI0_CLKI_posedge_posedge,
        HoldHigh       => thold_ADRI0_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C_FIFO",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_DATI0_CLKI_posedge ,
        TimingData     =>Tmkr_DATI0_CLKI_posedge  ,
        TestSignal     => DATI0_ipd,
        TestSignalName => "DATI0",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_DATI0_CLKI_posedge_posedge ,
        SetupLow       => tsetup_DATI0_CLKI_negedge_posedge,
        HoldLow        => thold_DATI0_CLKI_posedge_posedge,
        HoldHigh       => thold_DATI0_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C_FIFO",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_DATI1_CLKI_posedge ,
        TimingData     =>Tmkr_DATI1_CLKI_posedge  ,
        TestSignal     => DATI1_ipd,
        TestSignalName => "DATI1",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_DATI1_CLKI_posedge_posedge ,
        SetupLow       => tsetup_DATI1_CLKI_negedge_posedge,
        HoldLow        => thold_DATI1_CLKI_posedge_posedge,
        HoldHigh       => thold_DATI1_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C_FIFO",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_DATI2_CLKI_posedge ,
        TimingData     =>Tmkr_DATI2_CLKI_posedge  ,
        TestSignal     => DATI2_ipd,
        TestSignalName => "DATI2",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_DATI2_CLKI_posedge_posedge ,
        SetupLow       => tsetup_DATI2_CLKI_negedge_posedge,
        HoldLow        => thold_DATI2_CLKI_posedge_posedge,
        HoldHigh       => thold_DATI2_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C_FIFO",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_DATI3_CLKI_posedge ,
        TimingData     =>Tmkr_DATI3_CLKI_posedge  ,
        TestSignal     => DATI3_ipd,
        TestSignalName => "DATI3",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_DATI3_CLKI_posedge_posedge ,
        SetupLow       => tsetup_DATI3_CLKI_negedge_posedge,
        HoldLow        => thold_DATI3_CLKI_posedge_posedge,
        HoldHigh       => thold_DATI3_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C_FIFO",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_DATI4_CLKI_posedge ,
        TimingData     =>Tmkr_DATI4_CLKI_posedge  ,
        TestSignal     => DATI4_ipd,
        TestSignalName => "DATI4",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_DATI4_CLKI_posedge_posedge ,
        SetupLow       => tsetup_DATI4_CLKI_negedge_posedge,
        HoldLow        => thold_DATI4_CLKI_posedge_posedge,
        HoldHigh       => thold_DATI4_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C_FIFO",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_DATI5_CLKI_posedge ,
        TimingData     =>Tmkr_DATI5_CLKI_posedge  ,
        TestSignal     => DATI5_ipd,
        TestSignalName => "DATI5",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_DATI5_CLKI_posedge_posedge ,
        SetupLow       => tsetup_DATI5_CLKI_negedge_posedge,
        HoldLow        => thold_DATI5_CLKI_posedge_posedge,
        HoldHigh       => thold_DATI5_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C_FIFO",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_DATI6_CLKI_posedge ,
        TimingData     =>Tmkr_DATI6_CLKI_posedge  ,
        TestSignal     => DATI6_ipd,
        TestSignalName => "DATI6",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_DATI6_CLKI_posedge_posedge ,
        SetupLow       => tsetup_DATI6_CLKI_negedge_posedge,
        HoldLow        => thold_DATI6_CLKI_posedge_posedge,
        HoldHigh       => thold_DATI6_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C_FIFO",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_DATI7_CLKI_posedge ,
        TimingData     =>Tmkr_DATI7_CLKI_posedge  ,
        TestSignal     => DATI7_ipd,
        TestSignalName => "DATI7",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_DATI7_CLKI_posedge_posedge ,
        SetupLow       => tsetup_DATI7_CLKI_negedge_posedge,
        HoldLow        => thold_DATI7_CLKI_posedge_posedge,
        HoldHigh       => thold_DATI7_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C_FIFO",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_DATI8_CLKI_posedge ,
        TimingData     =>Tmkr_DATI8_CLKI_posedge  ,
        TestSignal     => DATI8_ipd,
        TestSignalName => "DATI8",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_DATI8_CLKI_posedge_posedge ,
        SetupLow       => tsetup_DATI8_CLKI_negedge_posedge,
        HoldLow        => thold_DATI8_CLKI_posedge_posedge,
        HoldHigh       => thold_DATI8_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C_FIFO",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_DATI9_CLKI_posedge ,
        TimingData     =>Tmkr_DATI9_CLKI_posedge  ,
        TestSignal     => DATI9_ipd,
        TestSignalName => "DATI9",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_DATI9_CLKI_posedge_posedge ,
        SetupLow       => tsetup_DATI9_CLKI_negedge_posedge,
        HoldLow        => thold_DATI9_CLKI_posedge_posedge,
        HoldHigh       => thold_DATI9_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C_FIFO",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_SCLI_CLKI_posedge ,
        TimingData     =>Tmkr_SCLI_CLKI_posedge  ,
        TestSignal     => SCLI_ipd,
        TestSignalName => "SCLI",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_SCLI_CLKI_posedge_posedge ,
        SetupLow       => tsetup_SCLI_CLKI_negedge_posedge,
        HoldLow        => thold_SCLI_CLKI_posedge_posedge,
        HoldHigh       => thold_SCLI_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_I2C_FIFO",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
 VitalPeriodPulseCheck (
        Violation      => Pviol_CLKI,
        PeriodData     => PInfo_CLKI,
        TestSignal     => CLKI_ipd,
        TestSignalName => "CLKI",
        TestDelay      => 0 ns,
        Period         => 0 ns,
        PulseWidthHigh => tpw_CLKI_posedge,
        PulseWidthLow  => tpw_CLKI_negedge,
        CheckEnabled   => true,
        HeaderMsg      => "/SB_I2C_FIFO",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
end if;
end process VITALBehavior;
VITALPathDelay   : process ( SCLO_sig, ACKO_sig, DATO0_sig, DATO1_sig, DATO2_sig, DATO3_sig, DATO4_sig, DATO5_sig, DATO6_sig, DATO7_sig, DATO8_sig, DATO9_sig, I2CIRQ_sig, I2CWKUP_sig, MRDCMPL_sig, RXFIFOAFULL_sig, RXFIFOEMPTY_sig, RXFIFOFULL_sig, SCLOE_sig, SDAO_sig, SDAOE_sig, SRWO_sig, TXFIFOAEMPTY_sig, TXFIFOEMPTY_sig, ADRI0_ipd, ADRI1_ipd, ADRI2_ipd, ADRI3_ipd, CLKI_ipd, CSI_ipd, DATI0_ipd, DATI1_ipd, DATI2_ipd, DATI3_ipd, DATI4_ipd, DATI5_ipd, DATI6_ipd, DATI7_ipd, DATI8_ipd, DATI9_ipd, FIFORST_ipd, SCLI_ipd, SDAI_ipd, STBI_ipd, WEI_ipd, TXFIFOFULL_sig)
variable SCLO_GlitchData : VitalGlitchDataType;
 variable SCLO_zd : std_logic :='X';
 variable ACKO_GlitchData : VitalGlitchDataType;
 variable ACKO_zd: std_logic :='X';
 variable DATO0_GlitchData : VitalGlitchDataType;
 variable DATO0_zd: std_logic :='X';
 variable DATO1_GlitchData : VitalGlitchDataType;
 variable DATO1_zd: std_logic :='X';
 variable DATO2_GlitchData : VitalGlitchDataType;
 variable DATO2_zd: std_logic :='X';
 variable DATO3_GlitchData : VitalGlitchDataType;
 variable DATO3_zd: std_logic :='X';
 variable DATO4_GlitchData : VitalGlitchDataType;
 variable DATO4_zd: std_logic :='X';
 variable DATO5_GlitchData : VitalGlitchDataType;
 variable DATO5_zd: std_logic :='X';
 variable DATO6_GlitchData : VitalGlitchDataType;
 variable DATO6_zd: std_logic :='X';
 variable DATO7_GlitchData : VitalGlitchDataType;
 variable DATO7_zd: std_logic :='X';
 variable DATO8_GlitchData : VitalGlitchDataType;
 variable DATO8_zd: std_logic :='X';
 variable DATO9_GlitchData : VitalGlitchDataType;
 variable DATO9_zd: std_logic :='X';
 variable I2CIRQ_GlitchData : VitalGlitchDataType;
 variable I2CIRQ_zd: std_logic :='X';
 variable I2CWKUP_GlitchData : VitalGlitchDataType;
 variable I2CWKUP_zd: std_logic :='X';
 variable MRDCMPL_GlitchData : VitalGlitchDataType;
 variable MRDCMPL_zd: std_logic :='X';
 variable RXFIFOAFULL_GlitchData : VitalGlitchDataType;
 variable RXFIFOAFULL_zd: std_logic :='X';
 variable RXFIFOEMPTY_GlitchData : VitalGlitchDataType;
 variable RXFIFOEMPTY_zd: std_logic :='X';
 variable RXFIFOFULL_GlitchData : VitalGlitchDataType;
 variable RXFIFOFULL_zd: std_logic :='X';
 variable SCLOE_GlitchData : VitalGlitchDataType;
 variable SCLOE_zd: std_logic :='X';
 variable SDAO_GlitchData : VitalGlitchDataType;
 variable SDAO_zd: std_logic :='X';
 variable SDAOE_GlitchData : VitalGlitchDataType;
 variable SDAOE_zd: std_logic :='X';
 variable SRWO_GlitchData : VitalGlitchDataType;
 variable SRWO_zd: std_logic :='X';
 variable TXFIFOAEMPTY_GlitchData : VitalGlitchDataType;
 variable TXFIFOAEMPTY_zd: std_logic :='X';
 variable TXFIFOEMPTY_GlitchData : VitalGlitchDataType;
 variable TXFIFOEMPTY_zd: std_logic :='X';
 variable TXFIFOFULL_GlitchData : VitalGlitchDataType;
 variable TXFIFOFULL_zd: std_logic :='X';
begin
SCLO_zd := SCLO_sig;
 ACKO_zd := ACKO_sig;
 DATO0_zd := DATO0_sig;
 DATO1_zd := DATO1_sig;
 DATO2_zd := DATO2_sig;
 DATO3_zd := DATO3_sig;
 DATO4_zd := DATO4_sig;
 DATO5_zd := DATO5_sig;
 DATO6_zd := DATO6_sig;
 DATO7_zd := DATO7_sig;
 DATO8_zd := DATO8_sig;
 DATO9_zd := DATO9_sig;
 I2CIRQ_zd := I2CIRQ_sig;
 I2CWKUP_zd := I2CWKUP_sig;
 MRDCMPL_zd := MRDCMPL_sig;
 SCLOE_zd := SCLOE_sig;
 SDAO_zd := SDAO_sig;
 SDAOE_zd := SDAOE_sig;
 SRWO_zd := SRWO_sig;
 RXFIFOAFULL_zd := RXFIFOAFULL_sig;
 RXFIFOEMPTY_zd := RXFIFOEMPTY_sig;
 RXFIFOFULL_zd := RXFIFOFULL_sig;
 TXFIFOAEMPTY_zd := TXFIFOAEMPTY_sig;
 TXFIFOEMPTY_zd := TXFIFOEMPTY_sig;
 TXFIFOFULL_zd := TXFIFOFULL_sig;

     VitalPathDelay01 (
	      OutSignal     => DATO0,
	      GlitchData    => DATO0_GlitchData,
	      OutSignalName => "DATO0",
	      OutTemp       => DATO0_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_DATO0_posedge, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => DATO1,
	      GlitchData    => DATO1_GlitchData,
	      OutSignalName => "DATO1",
	      OutTemp       => DATO1_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_DATO1_posedge, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => DATO2,
	      GlitchData    => DATO2_GlitchData,
	      OutSignalName => "DATO2",
	      OutTemp       => DATO2_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_DATO2_posedge, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => DATO3,
	      GlitchData    => DATO3_GlitchData,
	      OutSignalName => "DATO3",
	      OutTemp       => DATO3_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_DATO3_posedge, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => DATO4,
	      GlitchData    => DATO4_GlitchData,
	      OutSignalName => "DATO4",
	      OutTemp       => DATO4_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_DATO4_posedge, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => DATO5,
	      GlitchData    => DATO5_GlitchData,
	      OutSignalName => "DATO5",
	      OutTemp       => DATO5_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_DATO5_posedge, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => DATO6,
	      GlitchData    => DATO6_GlitchData,
	      OutSignalName => "DATO6",
	      OutTemp       => DATO6_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_DATO6_posedge, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => DATO7,
	      GlitchData    => DATO7_GlitchData,
	      OutSignalName => "DATO7",
	      OutTemp       => DATO7_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_DATO7_posedge, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => DATO8,
	      GlitchData    => DATO8_GlitchData,
	      OutSignalName => "DATO8",
	      OutTemp       => DATO8_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_DATO8_posedge, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => DATO9,
	      GlitchData    => DATO9_GlitchData,
	      OutSignalName => "DATO9",
	      OutTemp       => DATO9_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_DATO9_posedge, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => ACKO,
	      GlitchData    => ACKO_GlitchData,
	      OutSignalName => "ACKO",
	      OutTemp       => ACKO_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_ACKO_posedge, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => SRWO,
	      GlitchData    => SRWO_GlitchData,
	      OutSignalName => "SRWO",
	      OutTemp       => SRWO_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_SRWO_posedge, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => I2CIRQ,
	      GlitchData    => I2CIRQ_GlitchData,
	      OutSignalName => "I2CIRQ",
	      OutTemp       => I2CIRQ_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_I2CIRQ_posedge, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => I2CWKUP,
	      GlitchData    => I2CWKUP_GlitchData,
	      OutSignalName => "I2CWKUP",
	      OutTemp       => I2CWKUP_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_I2CWKUP_posedge, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => SCLO,
	      GlitchData    => SCLO_GlitchData,
	      OutSignalName => "SCLO",
	      OutTemp       => SCLO_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_SCLO_posedge, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => SCLOE,
	      GlitchData    => SCLOE_GlitchData,
	      OutSignalName => "SCLOE",
	      OutTemp       => SCLOE_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_SCLOE_posedge, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => SDAO,
	      GlitchData    => SDAO_GlitchData,
	      OutSignalName => "SDAO",
	      OutTemp       => SDAO_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_SDAO_posedge, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => SDAOE,
	      GlitchData    => SDAOE_GlitchData,
	      OutSignalName => "SDAOE",
	      OutTemp       => SDAOE_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_SDAOE_posedge, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
     
      VitalPathDelay01 (
	      OutSignal     => RXFIFOEMPTY,
	      GlitchData    => RXFIFOEMPTY_GlitchData,
	      OutSignalName => "RXFIFOEMPTY",
	      OutTemp       => RXFIFOEMPTY_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_RXFIFOEMPTY_posedge, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
     
      VitalPathDelay01 (
	      OutSignal     => RXFIFOAFULL,
	      GlitchData    => RXFIFOAFULL_GlitchData,
	      OutSignalName => "RXFIFOAFULL",
	      OutTemp       => RXFIFOAFULL_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_RXFIFOAFULL_posedge, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
     
      VitalPathDelay01 (
	      OutSignal     => RXFIFOFULL,
	      GlitchData    => RXFIFOFULL_GlitchData,
	      OutSignalName => "RXFIFOFULL",
	      OutTemp       => RXFIFOFULL_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_RXFIFOFULL_posedge, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
     
      VitalPathDelay01 (
	      OutSignal     => TXFIFOFULL,
	      GlitchData    => TXFIFOFULL_GlitchData,
	      OutSignalName => "TXFIFOFULL",
	      OutTemp       => TXFIFOFULL_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_TXFIFOFULL_posedge, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
     
      VitalPathDelay01 (
	      OutSignal     => TXFIFOAEMPTY,
	      GlitchData    => TXFIFOAEMPTY_GlitchData,
	      OutSignalName => "TXFIFOAEMPTY",
	      OutTemp       => TXFIFOAEMPTY_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_TXFIFOAEMPTY_posedge, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
     
       VitalPathDelay01 (
	      OutSignal     => TXFIFOEMPTY,
	      GlitchData    => TXFIFOEMPTY_GlitchData,
	      OutSignalName => "TXFIFOEMPTY",
	      OutTemp       => TXFIFOEMPTY_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_TXFIFOEMPTY_posedge, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

      VitalPathDelay01 (
	      OutSignal     => SDAO,
	      GlitchData    => SDAO_GlitchData,
	      OutSignalName => "SDAO",
	      OutTemp       => SDAO_zd,
	      Paths         => (0 => (SCLO_ipd'last_event, tpd_SCLO_SDAO_posedge, true),
                        1 => (SCLO_ipd'last_event, tpd_SCLO_SDAO_negedge, true),
						2 => (SCLI_ipd'last_event, tpd_SCLI_SDAO_negedge, true),
						3 => (SCLI_ipd'last_event, tpd_SCLI_SDAO_negedge, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => SDAOE,
	      GlitchData    => SDAOE_GlitchData,
	      OutSignalName => "SDAOE",
	      OutTemp       => SDAOE_zd,
	      Paths         => (0 => (SCLO_ipd'last_event, tpd_SCLO_SDAOE_posedge, true),
                        1 => (SCLO_ipd'last_event, tpd_SCLO_SDAOE_negedge, true),
						2 => (SCLI_ipd'last_event, tpd_SCLI_SDAOE_negedge, true),
						3 => (SCLI_ipd'last_event, tpd_SCLI_SDAOE_negedge, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
 end process VITALPathDelay;
end  SB_I2C_FIFO_V;		




-------------------------------------------------
---     	SB_IR_IP 		-------
------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;
use IEEE.VITAL_Timing.all; 
USE IEEE.numeric_std.ALL;
entity  SB_IR_IP  is
Generic 
(
    TimingChecksOn  : boolean := true;
    Xon   : boolean := true;					   
    MsgOn : boolean := false;
        tsetup_CSI_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       tsetup_CSI_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       thold_CSI_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       thold_CSI_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       tsetup_DENI_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       tsetup_DENI_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       thold_DENI_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       thold_DENI_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       tsetup_WEI_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       tsetup_WEI_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       thold_WEI_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       thold_WEI_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       tsetup_ADRI3_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       tsetup_ADRI3_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       thold_ADRI3_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       thold_ADRI3_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       tsetup_ADRI2_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       tsetup_ADRI2_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       thold_ADRI2_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       thold_ADRI2_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       tsetup_ADRI1_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       tsetup_ADRI1_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       thold_ADRI1_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       thold_ADRI1_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       tsetup_ADRI0_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       tsetup_ADRI0_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       thold_ADRI0_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       thold_ADRI0_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
	   tsetup_WDATA0_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       tsetup_WDATA0_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       thold_WDATA0_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       thold_WDATA0_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       tsetup_WDATA1_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       tsetup_WDATA1_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       thold_WDATA1_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       thold_WDATA1_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       tsetup_WDATA2_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       tsetup_WDATA2_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       thold_WDATA2_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       thold_WDATA2_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       tsetup_WDATA3_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       tsetup_WDATA3_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       thold_WDATA3_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       thold_WDATA3_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       tsetup_WDATA4_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       tsetup_WDATA4_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       thold_WDATA4_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       thold_WDATA4_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       tsetup_WDATA5_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       tsetup_WDATA5_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       thold_WDATA5_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       thold_WDATA5_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       tsetup_WDATA6_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       tsetup_WDATA6_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       thold_WDATA6_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       thold_WDATA6_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       tsetup_WDATA7_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       tsetup_WDATA7_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       thold_WDATA7_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       thold_WDATA7_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       tsetup_EXE_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       tsetup_EXE_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       thold_EXE_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       thold_EXE_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       tsetup_LEARN_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       tsetup_LEARN_CLKI_posedge_posedge : VitalDelayType:= 0 ns;
       thold_LEARN_CLKI_negedge_posedge : VitalDelayType := 0 ns;
       thold_LEARN_CLKI_posedge_posedge : VitalDelayType:= 0 ns;

        tpw_CLKI_posedge : VitalDelayType := 0 ns;
       tpw_CLKI_negedge : VitalDelayType := 0 ns;

        tpd_CLKI_BUSY : VitalDelayType01 := (0 ns, 0 ns);
       tpd_CLKI_BUSY_posedge : VitalDelayType01 := (0 ns, 0 ns);
       tpd_CLKI_DRDY : VitalDelayType01 := (0 ns, 0 ns);
       tpd_CLKI_DRDY_posedge : VitalDelayType01 := (0 ns, 0 ns);
       tpd_CLKI_ERR : VitalDelayType01 := (0 ns, 0 ns);
       tpd_CLKI_ERR_posedge : VitalDelayType01 := (0 ns, 0 ns);
       tpd_CLKI_IROUT : VitalDelayType01 := (0 ns, 0 ns);
       tpd_CLKI_IROUT_posedge : VitalDelayType01 := (0 ns, 0 ns);
       tpd_CLKI_RDATA0 : VitalDelayType01 := (0 ns, 0 ns);
       tpd_CLKI_RDATA0_posedge : VitalDelayType01 := (0 ns, 0 ns);
       tpd_CLKI_RDATA1 : VitalDelayType01 := (0 ns, 0 ns);
       tpd_CLKI_RDATA1_posedge : VitalDelayType01 := (0 ns, 0 ns);
       tpd_CLKI_RDATA2 : VitalDelayType01 := (0 ns, 0 ns);
       tpd_CLKI_RDATA2_posedge : VitalDelayType01 := (0 ns, 0 ns);
       tpd_CLKI_RDATA3 : VitalDelayType01 := (0 ns, 0 ns);
       tpd_CLKI_RDATA3_posedge : VitalDelayType01 := (0 ns, 0 ns);
       tpd_CLKI_RDATA4 : VitalDelayType01 := (0 ns, 0 ns);
       tpd_CLKI_RDATA4_posedge : VitalDelayType01 := (0 ns, 0 ns);
       tpd_CLKI_RDATA5 : VitalDelayType01 := (0 ns, 0 ns);
       tpd_CLKI_RDATA5_posedge : VitalDelayType01 := (0 ns, 0 ns);
       tpd_CLKI_RDATA6 : VitalDelayType01 := (0 ns, 0 ns);
       tpd_CLKI_RDATA6_posedge : VitalDelayType01 := (0 ns, 0 ns);
       tpd_CLKI_RDATA7 : VitalDelayType01 := (0 ns, 0 ns);
       tpd_CLKI_RDATA7_posedge : VitalDelayType01 := (0 ns, 0 ns);
  		tipd_ADRI0 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_ADRI1 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_ADRI2 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_ADRI3 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_CLKI 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_CSI 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_DENI 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_EXE 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_IRIN 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_LEARN 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_RST 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_WDATA0 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_WDATA1 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_WDATA2 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_WDATA3 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_WDATA4 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_WDATA5 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_WDATA6 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_WDATA7 	: VitalDelayType01 := (0.000 ns, 0.000 ns);
 		tipd_WEI 	: VitalDelayType01 := (0.000 ns, 0.000 ns)
);
port (
        ADRI0 : in std_logic;
		 ADRI1 : in std_logic;
		 ADRI2 : in std_logic;
		 ADRI3 : in std_logic;
		 CLKI : in std_logic;
		 CSI : in std_logic;
		 DENI : in std_logic;
		 EXE : in std_logic;
		 IRIN : in std_logic;
		 LEARN : in std_logic;
		 RST : in std_logic;
		 WDATA0 : in std_logic;
		 WDATA1 : in std_logic;
		 WDATA2 : in std_logic;
		 WDATA3 : in std_logic;
		 WDATA4 : in std_logic;
		 WDATA5 : in std_logic;
		 WDATA6 : in std_logic;
		 WDATA7 : in std_logic;
		 WEI : in std_logic;
        BUSY : out std_logic;
		 DRDY : out std_logic;
		 ERR : out std_logic;
		 IROUT : out std_logic;
		 RDATA0 : out std_logic;
		 RDATA1 : out std_logic;
		 RDATA2 : out std_logic;
		 RDATA3 : out std_logic;
		 RDATA4 : out std_logic;
		 RDATA5 : out std_logic;
		 RDATA6 : out std_logic;
		 RDATA7 : out std_logic
	);	 
attribute VITAL_LEVEL0 of
    SB_IR_IP  : entity is true;
end SB_IR_IP;

architecture SB_IR_IP_CORE_V of SB_IR_IP is
  attribute VITAL_LEVEL0 of
    SB_IR_IP_CORE_V: architecture is true;

          signal  ADRI0_ipd	: std_ulogic :='X' ;
       signal  ADRI1_ipd	: std_ulogic :='X' ;
       signal  ADRI2_ipd	: std_ulogic :='X' ;
       signal  ADRI3_ipd	: std_ulogic :='X' ;
       signal  CLKI_ipd	: std_ulogic :='X' ;
       signal  CSI_ipd	: std_ulogic :='X' ;
       signal  DENI_ipd	: std_ulogic :='X' ;
       signal  EXE_ipd	: std_ulogic :='X' ;
       signal  IRIN_ipd	: std_ulogic :='X' ;
       signal  LEARN_ipd	: std_ulogic :='X' ;
       signal  RST_ipd	: std_ulogic :='X' ;
       signal  WDATA0_ipd	: std_ulogic :='X' ;
       signal  WDATA1_ipd	: std_ulogic :='X' ;
       signal  WDATA2_ipd	: std_ulogic :='X' ;
       signal  WDATA3_ipd	: std_ulogic :='X' ;
       signal  WDATA4_ipd	: std_ulogic :='X' ;
       signal  WDATA5_ipd	: std_ulogic :='X' ;
       signal  WDATA6_ipd	: std_ulogic :='X' ;
       signal  WDATA7_ipd	: std_ulogic :='X' ;
       signal  WEI_ipd	: std_ulogic :='X' ;

      signal BUSY_sig: std_ulogic     := 'X';
        signal DRDY_sig: std_ulogic     := 'X';
        signal ERR_sig: std_ulogic     := 'X';
        signal IROUT_sig: std_ulogic     := 'X';
        signal RDATA0_sig: std_ulogic     := 'X';
        signal RDATA1_sig: std_ulogic     := 'X';
        signal RDATA2_sig: std_ulogic     := 'X';
        signal RDATA3_sig: std_ulogic     := 'X';
        signal RDATA4_sig: std_ulogic     := 'X';
        signal RDATA5_sig: std_ulogic     := 'X';
        signal RDATA6_sig: std_ulogic     := 'X';
        signal RDATA7_sig: std_ulogic     := 'X';
	component SB_IR_IP_CORE
		port ( ADRI0 : in std_logic;
		 ADRI1 : in std_logic;
		 ADRI2 : in std_logic;
		 ADRI3 : in std_logic;
		 CLKI : in std_logic;
		 CSI : in std_logic;
		 DENI : in std_logic;
		 EXE : in std_logic;
		 IRIN : in std_logic;
		 LEARN : in std_logic;
		 RST : in std_logic;
		 WDATA0 : in std_logic;
		 WDATA1 : in std_logic;
		 WDATA2 : in std_logic;
		 WDATA3 : in std_logic;
		 WDATA4 : in std_logic;
		 WDATA5 : in std_logic;
		 WDATA6 : in std_logic;
		 WDATA7 : in std_logic;
		 WEI : in std_logic;
       			 BUSY : out std_logic;
		 DRDY : out std_logic;
		 ERR : out std_logic;
		 IROUT : out std_logic;
		 RDATA0 : out std_logic;
		 RDATA1 : out std_logic;
		 RDATA2 : out std_logic;
		 RDATA3 : out std_logic;
		 RDATA4 : out std_logic;
		 RDATA5 : out std_logic;
		 RDATA6 : out std_logic;
		 RDATA7 : out std_logic
	                	);
	end component;

    begin
    WireDelay:block
    begin
      VitalWireDelay (ADRI0_ipd, ADRI0, tipd_ADRI0);
       VitalWireDelay (ADRI1_ipd, ADRI1, tipd_ADRI1);
       VitalWireDelay (ADRI2_ipd, ADRI2, tipd_ADRI2);
       VitalWireDelay (ADRI3_ipd, ADRI3, tipd_ADRI3);
       VitalWireDelay (CLKI_ipd, CLKI, tipd_CLKI);
       VitalWireDelay (CSI_ipd, CSI, tipd_CSI);
       VitalWireDelay (DENI_ipd, DENI, tipd_DENI);
       VitalWireDelay (EXE_ipd, EXE, tipd_EXE);
       VitalWireDelay (IRIN_ipd, IRIN, tipd_IRIN);
       VitalWireDelay (LEARN_ipd, LEARN, tipd_LEARN);
       VitalWireDelay (RST_ipd, RST, tipd_RST);
       VitalWireDelay (WDATA0_ipd, WDATA0, tipd_WDATA0);
       VitalWireDelay (WDATA1_ipd, WDATA1, tipd_WDATA1);
       VitalWireDelay (WDATA2_ipd, WDATA2, tipd_WDATA2);
       VitalWireDelay (WDATA3_ipd, WDATA3, tipd_WDATA3);
       VitalWireDelay (WDATA4_ipd, WDATA4, tipd_WDATA4);
       VitalWireDelay (WDATA5_ipd, WDATA5, tipd_WDATA5);
       VitalWireDelay (WDATA6_ipd, WDATA6, tipd_WDATA6);
       VitalWireDelay (WDATA7_ipd, WDATA7, tipd_WDATA7);
       VitalWireDelay (WEI_ipd, WEI, tipd_WEI);

    end block;
		INST: SB_IR_IP_CORE
		port map (
		 ADRI0 =>  ADRI0_ipd   ,
		  ADRI1 =>  ADRI1_ipd   ,
		  ADRI2 =>  ADRI2_ipd   ,
		  ADRI3 =>  ADRI3_ipd   ,
		  CLKI =>  CLKI_ipd   ,
		  CSI =>  CSI_ipd   ,
		  DENI =>  DENI_ipd   ,
		  EXE =>  EXE_ipd   ,
		  IRIN =>  IRIN_ipd   ,
		  LEARN =>  LEARN_ipd   ,
		  RST =>  RST_ipd   ,
		  WDATA0 =>  WDATA0_ipd   ,
		  WDATA1 =>  WDATA1_ipd   ,
		  WDATA2 =>  WDATA2_ipd   ,
		  WDATA3 =>  WDATA3_ipd   ,
		  WDATA4 =>  WDATA4_ipd   ,
		  WDATA5 =>  WDATA5_ipd   ,
		  WDATA6 =>  WDATA6_ipd   ,
		  WDATA7 =>  WDATA7_ipd   ,
		  WEI =>  WEI_ipd   ,
       	 	 BUSY =>  BUSY_sig   ,
		  DRDY =>  DRDY_sig   ,
		  ERR =>  ERR_sig   ,
		  IROUT =>  IROUT_sig   ,
		  RDATA0 =>  RDATA0_sig   ,
		  RDATA1 =>  RDATA1_sig   ,
		  RDATA2 =>  RDATA2_sig   ,
		  RDATA3 =>  RDATA3_sig   ,
		  RDATA4 =>  RDATA4_sig   ,
		  RDATA5 =>  RDATA5_sig   ,
		  RDATA6 =>  RDATA6_sig   ,
		  RDATA7 =>  RDATA7_sig   
		);
VITALBehavior   : process ( BUSY_sig, DRDY_sig, ERR_sig, IROUT_sig, RDATA0_sig, RDATA1_sig, RDATA2_sig, RDATA3_sig, RDATA4_sig, RDATA5_sig, RDATA6_sig, ADRI0_ipd, ADRI1_ipd, ADRI2_ipd, ADRI3_ipd, CLKI_ipd, CSI_ipd, DENI_ipd, EXE_ipd, IRIN_ipd, LEARN_ipd, RST_ipd, WDATA0_ipd,WDATA0_ipd, WDATA1_ipd, WDATA2_ipd, WDATA3_ipd, WDATA4_ipd, WDATA5_ipd, WDATA6_ipd, WDATA7_ipd, WEI_ipd, RDATA7_sig)

    variable      Tviol_CSI_CLKI_posedge : std_logic := '0';
     variable      Tmkr_CSI_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
     variable      Tviol_DENI_CLKI_posedge : std_logic := '0';
     variable      Tmkr_DENI_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
     variable      Tviol_WEI_CLKI_posedge : std_logic := '0';
     variable      Tmkr_WEI_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
     variable      Tviol_ADRI3_CLKI_posedge : std_logic := '0';
     variable      Tmkr_ADRI3_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
     variable      Tviol_ADRI2_CLKI_posedge : std_logic := '0';
     variable      Tmkr_ADRI2_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
     variable      Tviol_ADRI1_CLKI_posedge : std_logic := '0';
     variable      Tmkr_ADRI1_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
     variable      Tviol_ADRI0_CLKI_posedge : std_logic := '0';
     variable      Tmkr_ADRI0_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
	 variable      Tviol_WDATA0_CLKI_posedge : std_logic := '0';
     variable      Tmkr_WDATA0_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
     variable      Tviol_WDATA1_CLKI_posedge : std_logic := '0';
     variable      Tmkr_WDATA1_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
     variable      Tviol_WDATA2_CLKI_posedge : std_logic := '0';
     variable      Tmkr_WDATA2_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
     variable      Tviol_WDATA3_CLKI_posedge : std_logic := '0';
     variable      Tmkr_WDATA3_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
     variable      Tviol_WDATA4_CLKI_posedge : std_logic := '0';
     variable      Tmkr_WDATA4_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
     variable      Tviol_WDATA5_CLKI_posedge : std_logic := '0';
     variable      Tmkr_WDATA5_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
     variable      Tviol_WDATA6_CLKI_posedge : std_logic := '0';
     variable      Tmkr_WDATA6_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
     variable      Tviol_WDATA7_CLKI_posedge : std_logic := '0';
     variable      Tmkr_WDATA7_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
     variable      Tviol_EXE_CLKI_posedge : std_logic := '0';
     variable      Tmkr_EXE_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
     variable      Tviol_LEARN_CLKI_posedge : std_logic := '0';
     variable      Tmkr_LEARN_CLKI_posedge : VitalTimingDataType :=VitalTimingDataInit ;
 variable      Pviol_CLKI : std_logic := '0';
  variable      PInfo_CLKI : VitalPeriodDataType := VitalPeriodDataInit;
begin
if (TimingChecksOn) then
 VitalSetupHoldCheck (
        Violation      =>Tviol_CSI_CLKI_posedge ,
        TimingData     =>Tmkr_CSI_CLKI_posedge  ,
        TestSignal     => CSI_ipd,
        TestSignalName => "CSI",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_CSI_CLKI_posedge_posedge ,
        SetupLow       => tsetup_CSI_CLKI_negedge_posedge,
        HoldLow        => thold_CSI_CLKI_posedge_posedge,
        HoldHigh       => thold_CSI_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_IR_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_DENI_CLKI_posedge ,
        TimingData     =>Tmkr_DENI_CLKI_posedge  ,
        TestSignal     => DENI_ipd,
        TestSignalName => "DENI",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_DENI_CLKI_posedge_posedge ,
        SetupLow       => tsetup_DENI_CLKI_negedge_posedge,
        HoldLow        => thold_DENI_CLKI_posedge_posedge,
        HoldHigh       => thold_DENI_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_IR_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_WEI_CLKI_posedge ,
        TimingData     =>Tmkr_WEI_CLKI_posedge  ,
        TestSignal     => WEI_ipd,
        TestSignalName => "WEI",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WEI_CLKI_posedge_posedge ,
        SetupLow       => tsetup_WEI_CLKI_negedge_posedge,
        HoldLow        => thold_WEI_CLKI_posedge_posedge,
        HoldHigh       => thold_WEI_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_IR_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_ADRI3_CLKI_posedge ,
        TimingData     =>Tmkr_ADRI3_CLKI_posedge  ,
        TestSignal     => ADRI3_ipd,
        TestSignalName => "ADRI3",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_ADRI3_CLKI_posedge_posedge ,
        SetupLow       => tsetup_ADRI3_CLKI_negedge_posedge,
        HoldLow        => thold_ADRI3_CLKI_posedge_posedge,
        HoldHigh       => thold_ADRI3_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_IR_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_ADRI2_CLKI_posedge ,
        TimingData     =>Tmkr_ADRI2_CLKI_posedge  ,
        TestSignal     => ADRI2_ipd,
        TestSignalName => "ADRI2",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_ADRI2_CLKI_posedge_posedge ,
        SetupLow       => tsetup_ADRI2_CLKI_negedge_posedge,
        HoldLow        => thold_ADRI2_CLKI_posedge_posedge,
        HoldHigh       => thold_ADRI2_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_IR_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_ADRI1_CLKI_posedge ,
        TimingData     =>Tmkr_ADRI1_CLKI_posedge  ,
        TestSignal     => ADRI1_ipd,
        TestSignalName => "ADRI1",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_ADRI1_CLKI_posedge_posedge ,
        SetupLow       => tsetup_ADRI1_CLKI_negedge_posedge,
        HoldLow        => thold_ADRI1_CLKI_posedge_posedge,
        HoldHigh       => thold_ADRI1_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_IR_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_ADRI0_CLKI_posedge ,
        TimingData     =>Tmkr_ADRI0_CLKI_posedge  ,
        TestSignal     => ADRI0_ipd,
        TestSignalName => "ADRI0",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_ADRI0_CLKI_posedge_posedge ,
        SetupLow       => tsetup_ADRI0_CLKI_negedge_posedge,
        HoldLow        => thold_ADRI0_CLKI_posedge_posedge,
        HoldHigh       => thold_ADRI0_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_IR_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
	VitalSetupHoldCheck (
        Violation      =>Tviol_WDATA0_CLKI_posedge ,
        TimingData     =>Tmkr_WDATA0_CLKI_posedge  ,
        TestSignal     => WDATA0_ipd,
        TestSignalName => "WDATA0",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA0_CLKI_posedge_posedge ,
        SetupLow       => tsetup_WDATA0_CLKI_negedge_posedge,
        HoldLow        => thold_WDATA0_CLKI_posedge_posedge,
        HoldHigh       => thold_WDATA0_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_IR_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_WDATA1_CLKI_posedge ,
        TimingData     =>Tmkr_WDATA1_CLKI_posedge  ,
        TestSignal     => WDATA1_ipd,
        TestSignalName => "WDATA1",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA1_CLKI_posedge_posedge ,
        SetupLow       => tsetup_WDATA1_CLKI_negedge_posedge,
        HoldLow        => thold_WDATA1_CLKI_posedge_posedge,
        HoldHigh       => thold_WDATA1_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_IR_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_WDATA2_CLKI_posedge ,
        TimingData     =>Tmkr_WDATA2_CLKI_posedge  ,
        TestSignal     => WDATA2_ipd,
        TestSignalName => "WDATA2",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA2_CLKI_posedge_posedge ,
        SetupLow       => tsetup_WDATA2_CLKI_negedge_posedge,
        HoldLow        => thold_WDATA2_CLKI_posedge_posedge,
        HoldHigh       => thold_WDATA2_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_IR_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_WDATA3_CLKI_posedge ,
        TimingData     =>Tmkr_WDATA3_CLKI_posedge  ,
        TestSignal     => WDATA3_ipd,
        TestSignalName => "WDATA3",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA3_CLKI_posedge_posedge ,
        SetupLow       => tsetup_WDATA3_CLKI_negedge_posedge,
        HoldLow        => thold_WDATA3_CLKI_posedge_posedge,
        HoldHigh       => thold_WDATA3_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_IR_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_WDATA4_CLKI_posedge ,
        TimingData     =>Tmkr_WDATA4_CLKI_posedge  ,
        TestSignal     => WDATA4_ipd,
        TestSignalName => "WDATA4",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA4_CLKI_posedge_posedge ,
        SetupLow       => tsetup_WDATA4_CLKI_negedge_posedge,
        HoldLow        => thold_WDATA4_CLKI_posedge_posedge,
        HoldHigh       => thold_WDATA4_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_IR_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_WDATA5_CLKI_posedge ,
        TimingData     =>Tmkr_WDATA5_CLKI_posedge  ,
        TestSignal     => WDATA5_ipd,
        TestSignalName => "WDATA5",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA5_CLKI_posedge_posedge ,
        SetupLow       => tsetup_WDATA5_CLKI_negedge_posedge,
        HoldLow        => thold_WDATA5_CLKI_posedge_posedge,
        HoldHigh       => thold_WDATA5_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_IR_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_WDATA6_CLKI_posedge ,
        TimingData     =>Tmkr_WDATA6_CLKI_posedge  ,
        TestSignal     => WDATA6_ipd,
        TestSignalName => "WDATA6",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA6_CLKI_posedge_posedge ,
        SetupLow       => tsetup_WDATA6_CLKI_negedge_posedge,
        HoldLow        => thold_WDATA6_CLKI_posedge_posedge,
        HoldHigh       => thold_WDATA6_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_IR_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_WDATA7_CLKI_posedge ,
        TimingData     =>Tmkr_WDATA7_CLKI_posedge  ,
        TestSignal     => WDATA7_ipd,
        TestSignalName => "WDATA7",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_WDATA7_CLKI_posedge_posedge ,
        SetupLow       => tsetup_WDATA7_CLKI_negedge_posedge,
        HoldLow        => thold_WDATA7_CLKI_posedge_posedge,
        HoldHigh       => thold_WDATA7_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_IR_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_EXE_CLKI_posedge ,
        TimingData     =>Tmkr_EXE_CLKI_posedge  ,
        TestSignal     => EXE_ipd,
        TestSignalName => "EXE",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_EXE_CLKI_posedge_posedge ,
        SetupLow       => tsetup_EXE_CLKI_negedge_posedge,
        HoldLow        => thold_EXE_CLKI_posedge_posedge,
        HoldHigh       => thold_EXE_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_IR_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
  VitalSetupHoldCheck (
        Violation      =>Tviol_LEARN_CLKI_posedge ,
        TimingData     =>Tmkr_LEARN_CLKI_posedge  ,
        TestSignal     => LEARN_ipd,
        TestSignalName => "LEARN",
        TestDelay      => 0 ns,
        RefSignal      => CLKI_ipd,
        RefSignalName  => "CLKI",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_LEARN_CLKI_posedge_posedge ,
        SetupLow       => tsetup_LEARN_CLKI_negedge_posedge,
        HoldLow        => thold_LEARN_CLKI_posedge_posedge,
        HoldHigh       => thold_LEARN_CLKI_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_IR_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
 VitalPeriodPulseCheck (
        Violation      => Pviol_CLKI,
        PeriodData     => PInfo_CLKI,
        TestSignal     => CLKI_ipd,
        TestSignalName => "CLKI",
        TestDelay      => 0 ns,
        Period         => 0 ns,
        PulseWidthHigh => tpw_CLKI_posedge,
        PulseWidthLow  => tpw_CLKI_negedge,
        CheckEnabled   => true,
        HeaderMsg      => "/SB_IR_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);
end if;
end process VITALBehavior;
VITALPathDelay   : process ( BUSY_sig, DRDY_sig, ERR_sig, IROUT_sig, RDATA0_sig, RDATA1_sig, RDATA2_sig, RDATA3_sig, RDATA4_sig, RDATA5_sig, RDATA6_sig, ADRI0_ipd, ADRI1_ipd, ADRI2_ipd, ADRI3_ipd, CLKI_ipd, CSI_ipd, DENI_ipd, EXE_ipd, IRIN_ipd, LEARN_ipd, RST_ipd, WDATA0_ipd, WDATA1_ipd, WDATA2_ipd, WDATA3_ipd, WDATA4_ipd, WDATA5_ipd, WDATA6_ipd, WDATA7_ipd, WEI_ipd, RDATA7_sig)
variable BUSY_GlitchData : VitalGlitchDataType;
 variable BUSY_zd: std_logic :='X';
 variable DRDY_GlitchData : VitalGlitchDataType;
 variable DRDY_zd: std_logic :='X';
 variable ERR_GlitchData : VitalGlitchDataType;
 variable ERR_zd: std_logic :='X';
 variable IROUT_GlitchData : VitalGlitchDataType;
 variable IROUT_zd: std_logic :='X';
 variable RDATA0_GlitchData : VitalGlitchDataType;
 variable RDATA0_zd: std_logic :='X';
 variable RDATA1_GlitchData : VitalGlitchDataType;
 variable RDATA1_zd: std_logic :='X';
 variable RDATA2_GlitchData : VitalGlitchDataType;
 variable RDATA2_zd: std_logic :='X';
 variable RDATA3_GlitchData : VitalGlitchDataType;
 variable RDATA3_zd: std_logic :='X';
 variable RDATA4_GlitchData : VitalGlitchDataType;
 variable RDATA4_zd: std_logic :='X';
 variable RDATA5_GlitchData : VitalGlitchDataType;
 variable RDATA5_zd: std_logic :='X';
 variable RDATA6_GlitchData : VitalGlitchDataType;
 variable RDATA6_zd: std_logic :='X';
 variable RDATA7_GlitchData : VitalGlitchDataType;
 variable RDATA7_zd: std_logic :='X';
begin
BUSY_zd := BUSY_sig;
 DRDY_zd := DRDY_sig;
 ERR_zd := ERR_sig;
 IROUT_zd := IROUT_sig;
 RDATA0_zd := RDATA0_sig;
 RDATA1_zd := RDATA1_sig;
 RDATA2_zd := RDATA2_sig;
 RDATA3_zd := RDATA3_sig;
 RDATA4_zd := RDATA4_sig;
 RDATA5_zd := RDATA5_sig;
 RDATA6_zd := RDATA6_sig;
 RDATA7_zd := RDATA7_sig;

     VitalPathDelay01 (
	      OutSignal     => RDATA0,
	      GlitchData    => RDATA0_GlitchData,
	      OutSignalName => "RDATA0",
	      OutTemp       => RDATA0_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_RDATA0, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => RDATA1,
	      GlitchData    => RDATA1_GlitchData,
	      OutSignalName => "RDATA1",
	      OutTemp       => RDATA1_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_RDATA1, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => RDATA2,
	      GlitchData    => RDATA2_GlitchData,
	      OutSignalName => "RDATA2",
	      OutTemp       => RDATA2_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_RDATA2, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => RDATA3,
	      GlitchData    => RDATA3_GlitchData,
	      OutSignalName => "RDATA3",
	      OutTemp       => RDATA3_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_RDATA3, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => RDATA4,
	      GlitchData    => RDATA4_GlitchData,
	      OutSignalName => "RDATA4",
	      OutTemp       => RDATA4_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_RDATA4, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => RDATA5,
	      GlitchData    => RDATA5_GlitchData,
	      OutSignalName => "RDATA5",
	      OutTemp       => RDATA5_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_RDATA5, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => RDATA6,
	      GlitchData    => RDATA6_GlitchData,
	      OutSignalName => "RDATA6",
	      OutTemp       => RDATA6_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_RDATA6, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => RDATA7,
	      GlitchData    => RDATA7_GlitchData,
	      OutSignalName => "RDATA7",
	      OutTemp       => RDATA7_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_RDATA7, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => BUSY,
	      GlitchData    => BUSY_GlitchData,
	      OutSignalName => "BUSY",
	      OutTemp       => BUSY_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_BUSY, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => DRDY,
	      GlitchData    => DRDY_GlitchData,
	      OutSignalName => "DRDY",
	      OutTemp       => DRDY_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_DRDY, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => ERR,
	      GlitchData    => ERR_GlitchData,
	      OutSignalName => "ERR",
	      OutTemp       => ERR_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_ERR, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
      VitalPathDelay01 (
	      OutSignal     => IROUT,
	      GlitchData    => IROUT_GlitchData,
	      OutSignalName => "IROUT",
	      OutTemp       => IROUT_zd,
	      Paths         => (0 => (CLKI_ipd'last_event, tpd_CLKI_IROUT, true)
),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);
 end process VITALPathDelay;
end  SB_IR_IP_CORE_V;		



-------------------------------------------------
---     	SB_RGB_IP 		-------
-----------------------------------------------

library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use work.std_logic_SBT.all;
entity  SB_RGB_IP  is
port (
CLK: in std_logic;
RST: in std_logic;
PARAMSOK: in std_logic;
RGBCOLOR: in std_logic_vector (3 downto 0); 
BRIGHTNESS: in std_logic_vector (3 downto 0); 
BREATHRAMP: in std_logic_vector (3 downto 0); 
BLINKRATE: in std_logic_vector (3 downto 0); 
REDPWM: out std_logic;
GREENPWM:out std_logic;
BLUEPWM:out std_logic
  ); 
end SB_RGB_IP;

architecture Behavior_SB_RGB_IP of SB_RGB_IP is

	component LED_control
		port ( 
		clk27M: in std_logic;
		rst: in std_logic;
		params_ok: in std_logic;
		RGB_color: in std_logic_vector (3 downto 0); 
		Brightness: in std_logic_vector (3 downto 0); 
		BreatheRamp: in std_logic_vector (3 downto 0); 
		BlinkRate: in std_logic_vector (3 downto 0); 
		red_pwm: out std_logic;
		grn_pwm:out std_logic;
		blu_pwm:out std_logic
	                	);
	end component;
	begin
		INST: LED_control
		port map (
		 clk27M =>  CLK   ,
		  params_ok =>  PARAMSOK   ,
		  rst =>  RST   ,
		  RGB_color =>RGBCOLOR,
		  Brightness =>BRIGHTNESS,
		  BlinkRate =>BLINKRATE,
		  BreatheRamp=>BREATHRAMP,
       	 	 blu_pwm =>  BLUEPWM   ,
		  grn_pwm =>  GREENPWM   ,
		  red_pwm =>  REDPWM   
		);
end  Behavior_SB_RGB_IP;		
--------------------------------------------------
---     	SB_LEDDA_IP 		-------
------------------------------------------------

library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use IEEE.VITAL_Primitives.all;
use IEEE.VITAL_Timing.all;
use work.std_logic_SBT.all;
entity  SB_LEDDA_IP  is 

generic (
	TimingChecksOn  	: boolean := true;
	Xon   			: boolean := true;
	MsgOn 			: boolean := true;

	tipd_LEDDCS:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDCLK:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDDAT7:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDDAT6:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDDAT5:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDDAT4:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDDAT3:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDDAT2:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDDAT1:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDDAT0:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDADDR3:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDADDR2:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDADDR1:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDADDR0:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDDEN:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDEXE:VitalDelayType01 := (0 ns, 0 ns);
	tipd_LEDDRST:VitalDelayType01 := (0 ns, 0 ns);
	tpd_LEDDCLK_LEDDON_posedge :VitalDelayType01 := (100 ns, 100 ns);
	tpd_LEDDCLK_PWMOUT0_posedge :VitalDelayType01 := (100 ns, 100 ns);
	tpd_LEDDCLK_PWMOUT1_posedge :VitalDelayType01 := (100 ns, 100 ns);
	tpd_LEDDCLK_PWMOUT2_posedge :VitalDelayType01 := (100 ns, 100 ns);
	
	tsetup_LEDDCS_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;	
	tsetup_LEDDCS_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDEN_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;	
	tsetup_LEDDDEN_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDEXE_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;	
	tsetup_LEDDEXE_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDADDR0_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDADDR0_LEDDCLK_negedge_posedge :VitalDelayType := 0 ns;
	tsetup_LEDDADDR1_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDADDR1_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDADDR2_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDADDR2_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDADDR3_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDADDR3_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	
	tsetup_LEDDDAT0_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDAT0_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDAT1_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDAT1_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDAT2_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDAT2_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDAT3_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDAT3_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDAT4_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDAT4_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDAT5_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDAT5_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDAT6_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDAT6_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDAT7_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	tsetup_LEDDDAT7_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	
	thold_LEDDCS_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;	
	thold_LEDDCS_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDEN_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;	
	thold_LEDDDEN_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDEXE_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;	
	thold_LEDDEXE_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDADDR0_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDADDR0_LEDDCLK_negedge_posedge :VitalDelayType := 0 ns;
	thold_LEDDADDR1_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDADDR1_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDADDR2_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDADDR2_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDADDR3_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDADDR3_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	
	thold_LEDDDAT0_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDAT0_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDAT1_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDAT1_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDAT2_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDAT2_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDAT3_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDAT3_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDAT4_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDAT4_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDAT5_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDAT5_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDAT6_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDAT6_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDAT7_LEDDCLK_posedge_posedge : VitalDelayType := 0 ns;
	thold_LEDDDAT7_LEDDCLK_negedge_posedge : VitalDelayType := 0 ns
	
);
 
port(
	PWMOUT0 : out std_logic;	
	PWMOUT1 : out std_logic;
	PWMOUT2 : out std_logic;
	LEDDON : out std_logic; 
	LEDDCS:in std_logic;
	LEDDCLK:in std_logic;
	LEDDDAT7:in std_logic;
	LEDDDAT6:in std_logic;
	LEDDDAT5:in std_logic;
	LEDDDAT4:in std_logic;
	LEDDDAT3:in std_logic;
	LEDDDAT2:in std_logic;
	LEDDDAT1:in std_logic;
	LEDDDAT0:in std_logic;
	LEDDADDR3:in std_logic;
	LEDDADDR2:in std_logic;
	LEDDADDR1:in std_logic;
	LEDDADDR0:in std_logic;
	LEDDDEN:in std_logic;
	LEDDEXE:in std_logic;
	LEDDRST:in std_logic
    );
	attribute VITAL_LEVEL0 of			    
    SB_LEDDA_IP  : entity is true;
end SB_LEDDA_IP ;

architecture SB_LEDDA_IP_V of SB_LEDDA_IP is
attribute VITAL_LEVEL0 of
    SB_LEDDA_IP_V : architecture is true;

SIGNAL LEDD_ADDR: std_logic_vector (3 downto 0);   
SIGNAL LEDD_DAT: std_logic_vector (7 downto 0);

	signal  PWMOUT0_sig  : std_ulogic	:='X';	
	signal  PWMOUT1_sig  : std_ulogic	:='X';
	signal  PWMOUT2_sig  : std_ulogic	:='X';
	signal  LEDDON_sig  : std_ulogic	:='X'; 
	
	signal  LEDDCS_ipd: std_ulogic := 'X';
	signal  LEDDCLK_ipd: std_ulogic := 'X';
	signal  LEDDDAT7_ipd: std_ulogic := 'X';
	signal  LEDDDAT6_ipd: std_ulogic := 'X';
	signal  LEDDDAT5_ipd: std_ulogic := 'X';
	signal  LEDDDAT4_ipd: std_ulogic := 'X';
	signal  LEDDDAT3_ipd: std_ulogic := 'X';
	signal  LEDDDAT2_ipd: std_ulogic := 'X';
	signal  LEDDDAT1_ipd: std_ulogic := 'X';
	signal  LEDDDAT0_ipd: std_ulogic := 'X';
	signal  LEDDADDR3_ipd: std_ulogic := 'X';
	signal  LEDDADDR2_ipd: std_ulogic := 'X';
	signal  LEDDADDR1_ipd: std_ulogic := 'X';
	signal  LEDDADDR0_ipd: std_ulogic := 'X';
	signal  LEDDDEN_ipd: std_ulogic := 'X';
	signal  LEDDEXE_ipd: std_ulogic := 'X';
	signal  LEDDRST_ipd: std_ulogic := 'X';
	signal ledd_rst:std_logic :='1';

component ledd_ip 
port	(
	pwm_out_r:out std_logic;
	pwm_out_g:out std_logic;
	pwm_out_b:out std_logic; 
	ledd_on :out std_logic;
	ledd_rst_async :in std_logic; 
	ledd_clk :in std_logic;
	ledd_cs :in std_logic;
	ledd_den :in std_logic; 
	ledd_adr :in std_logic_vector (3 downto 0); 
	ledd_dat :in std_logic_vector (7 downto 0);
    ledd_exe :in std_logic
   );
end component;

begin
	-- reset irip for 100ns -- 
process
begin
	wait for 100ns;
	ledd_rst <= '0';
	wait; 	
end process;

WireDelay : block
  begin
    VitalWireDelay (LEDDCS_ipd, LEDDCS, tipd_LEDDCS);
	VitalWireDelay (LEDDCLK_ipd, LEDDCLK, tipd_LEDDCLK);
	VitalWireDelay (LEDDDAT7_ipd, LEDDDAT7, tipd_LEDDDAT7);
	VitalWireDelay (LEDDDAT6_ipd, LEDDDAT6, tipd_LEDDDAT6);
	VitalWireDelay (LEDDDAT5_ipd, LEDDDAT5, tipd_LEDDDAT5);
	VitalWireDelay (LEDDDAT4_ipd, LEDDDAT4, tipd_LEDDDAT4);
	VitalWireDelay (LEDDDAT3_ipd, LEDDDAT3, tipd_LEDDDAT3);
	VitalWireDelay (LEDDDAT2_ipd, LEDDDAT2, tipd_LEDDDAT2);
	VitalWireDelay (LEDDDAT1_ipd, LEDDDAT1, tipd_LEDDDAT1);
	VitalWireDelay (LEDDDAT0_ipd, LEDDDAT0, tipd_LEDDDAT0);
	VitalWireDelay (LEDDADDR3_ipd, LEDDADDR3, tipd_LEDDADDR3);
	VitalWireDelay (LEDDADDR2_ipd, LEDDADDR2, tipd_LEDDADDR2);
	VitalWireDelay (LEDDADDR1_ipd, LEDDADDR1, tipd_LEDDADDR1);
	VitalWireDelay (LEDDADDR0_ipd, LEDDADDR0, tipd_LEDDADDR0);
	VitalWireDelay (LEDDDEN_ipd, LEDDDEN, tipd_LEDDDEN);
	VitalWireDelay (LEDDEXE_ipd, LEDDEXE, tipd_LEDDEXE);
	VitalWireDelay (LEDDRST_ipd, LEDDRST, tipd_LEDDRST);
	
  end block;

LS: ledd_ip 
port map(
	pwm_out_r =>PWMOUT0_sig  ,
	pwm_out_g =>PWMOUT1_sig  ,
	pwm_out_b =>PWMOUT2_sig  , 
	ledd_on  =>LEDDON_sig  ,
	ledd_rst_async  =>ledd_rst  , 
	ledd_clk  => LEDDCLK_ipd ,
	ledd_cs  => LEDDCS_ipd ,
	ledd_den  => LEDDDEN_ipd , 
	ledd_adr =>LEDD_ADDR,    
	ledd_dat  =>LEDD_DAT,    
    ledd_exe => LEDDEXE_ipd   
);
LEDD_ADDR<=(LEDDADDR3_ipd,LEDDADDR2_ipd,LEDDADDR1_ipd,LEDDADDR0_ipd) ; 
LEDD_DAT<=(LEDDDAT7_ipd,LEDDDAT6_ipd,LEDDDAT5_ipd,LEDDDAT4_ipd,LEDDDAT3_ipd,LEDDDAT2_ipd,LEDDDAT1_ipd,LEDDDAT0_ipd);

VITALBehavior : process(  PWMOUT0_sig,PWMOUT1_sig, PWMOUT2_sig,LEDDON_sig,LEDDCS_ipd,LEDDCLK_ipd,LEDDDAT7_ipd,LEDDDAT6_ipd,
	  LEDDDAT5_ipd,LEDDDAT4_ipd,LEDDDAT3_ipd,LEDDDAT2_ipd,LEDDDAT1_ipd,LEDDDAT0_ipd,LEDDADDR3_ipd,LEDDADDR2_ipd,LEDDADDR1_ipd,
	  LEDDADDR0_ipd,LEDDDEN_ipd,LEDDEXE_ipd,LEDDRST_ipd)

	variable Tviol_LEDDCS_LEDDCLK_posedge : std_logic := '0';	
	variable Tviol_LEDDDEN_LEDDCLK_posedge : std_logic := '0';	
	variable Tviol_LEDDEXE_LEDDCLK_posedge : std_logic := '0';	
	variable Tviol_LEDDADDR0_LEDDCLK_posedge : std_logic := '0';
	variable Tviol_LEDDADDR1_LEDDCLK_posedge : std_logic := '0';
	variable Tviol_LEDDADDR2_LEDDCLK_posedge : std_logic := '0';
	variable Tviol_LEDDADDR3_LEDDCLK_posedge : std_logic := '0';

	variable Tviol_LEDDDAT0_LEDDCLK_posedge : std_logic := '0';
	variable Tviol_LEDDDAT1_LEDDCLK_posedge : std_logic := '0';
	variable Tviol_LEDDDAT2_LEDDCLK_posedge : std_logic := '0';
	variable Tviol_LEDDDAT3_LEDDCLK_posedge : std_logic := '0';
	variable Tviol_LEDDDAT4_LEDDCLK_posedge : std_logic := '0';
	variable Tviol_LEDDDAT5_LEDDCLK_posedge : std_logic := '0';
	variable Tviol_LEDDDAT6_LEDDCLK_posedge : std_logic := '0';
	variable Tviol_LEDDDAT7_LEDDCLK_posedge : std_logic := '0';
	
	variable Tmkr_LEDDCS_LEDDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;	
	variable Tmkr_LEDDDEN_LEDDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;	
	variable Tmkr_LEDDEXE_LEDDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;	
	variable Tmkr_LEDDADDR0_LEDDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LEDDADDR1_LEDDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LEDDADDR2_LEDDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LEDDADDR3_LEDDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;

	variable Tmkr_LEDDDAT0_LEDDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LEDDDAT1_LEDDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LEDDDAT2_LEDDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LEDDDAT3_LEDDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LEDDDAT4_LEDDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LEDDDAT5_LEDDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LEDDDAT6_LEDDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LEDDDAT7_LEDDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable LEDDON_GlitchData : VitalGlitchDataType;  
	variable PWMOUT0_GlitchData : VitalGlitchDataType;
	variable PWMOUT1_GlitchData : VitalGlitchDataType;
	variable PWMOUT2_GlitchData : VitalGlitchDataType;				 
	variable PWMOUT0_zd :std_ulogic :='X';
	variable PWMOUT1_zd :std_ulogic :='X';
	variable PWMOUT2_zd :std_ulogic :='X'; 
	variable LEDDON_zd : std_ulogic :='X';

begin	  	
	PWMOUT0_zd:=PWMOUT0_sig;
	PWMOUT1_zd:=PWMOUT1_sig;
	PWMOUT2_zd:=PWMOUT2_sig;
	LEDDON_zd :=LEDDON_sig;
	if (TimingChecksOn) then
      VitalSetupHoldCheck (
        Violation      => Tviol_LEDDCS_LEDDCLK_posedge,
        TimingData     => Tmkr_LEDDCS_LEDDCLK_posedge,
        TestSignal     => LEDDCS_ipd,
        TestSignalName => "LEDDCS",
        TestDelay      => 0 ns,
        RefSignal      => LEDDCLK_ipd,
        RefSignalName  => "LEDDCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_LEDDCS_LEDDCLK_posedge_posedge,
        SetupLow       => tsetup_LEDDCS_LEDDCLK_negedge_posedge,
        HoldLow        => thold_LEDDCS_LEDDCLK_posedge_posedge,
        HoldHigh       => thold_LEDDCS_LEDDCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_LEDDA_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	  
	      VitalSetupHoldCheck (
        Violation      => Tviol_LEDDDEN_LEDDCLK_posedge,
        TimingData     => Tmkr_LEDDDEN_LEDDCLK_posedge,
        TestSignal     => LEDDDEN_ipd,
        TestSignalName => "LEDDDEN",
        TestDelay      => 0 ns,
        RefSignal      => LEDDCLK_ipd,
        RefSignalName  => "LEDDCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_LEDDDEN_LEDDCLK_posedge_posedge,
        SetupLow       => tsetup_LEDDDEN_LEDDCLK_negedge_posedge,
        HoldLow        => thold_LEDDDEN_LEDDCLK_posedge_posedge,
        HoldHigh       => thold_LEDDDEN_LEDDCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_LEDDA_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	 
		
		      VitalSetupHoldCheck (
        Violation      => Tviol_LEDDEXE_LEDDCLK_posedge,
        TimingData     => Tmkr_LEDDEXE_LEDDCLK_posedge,
        TestSignal     => LEDDEXE_ipd,
        TestSignalName => "LEDDEXE",
        TestDelay      => 0 ns,
        RefSignal      => LEDDCLK_ipd,
        RefSignalName  => "LEDDCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_LEDDEXE_LEDDCLK_posedge_posedge,
        SetupLow       => tsetup_LEDDEXE_LEDDCLK_negedge_posedge,
        HoldLow        => thold_LEDDEXE_LEDDCLK_posedge_posedge,
        HoldHigh       => thold_LEDDEXE_LEDDCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_LEDDA_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	 
		
		      VitalSetupHoldCheck (
        Violation      => Tviol_LEDDADDR0_LEDDCLK_posedge,
        TimingData     => Tmkr_LEDDADDR0_LEDDCLK_posedge,
        TestSignal     => LEDDADDR0_ipd,	 
        TestSignalName => "LEDDADDR0",
        TestDelay      => 0 ns,
        RefSignal      => LEDDCLK_ipd,
        RefSignalName  => "LEDDCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_LEDDADDR0_LEDDCLK_posedge_posedge,
        SetupLow       => tsetup_LEDDADDR0_LEDDCLK_negedge_posedge,
        HoldLow        => thold_LEDDADDR0_LEDDCLK_posedge_posedge,
        HoldHigh       => thold_LEDDADDR0_LEDDCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_LEDDA_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	 
		
		      VitalSetupHoldCheck (
        Violation      => Tviol_LEDDADDR1_LEDDCLK_posedge,
        TimingData     => Tmkr_LEDDADDR1_LEDDCLK_posedge,
        TestSignal     => LEDDADDR1_ipd,
        TestSignalName => "LEDDADDR1",
        TestDelay      => 0 ns,
        RefSignal      => LEDDCLK_ipd,
        RefSignalName  => "LEDDCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_LEDDADDR1_LEDDCLK_posedge_posedge,
        SetupLow       => tsetup_LEDDADDR1_LEDDCLK_negedge_posedge,
        HoldLow        => thold_LEDDADDR1_LEDDCLK_posedge_posedge,
        HoldHigh       => thold_LEDDADDR1_LEDDCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_LEDDA_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
		
		      VitalSetupHoldCheck (
        Violation      => Tviol_LEDDADDR2_LEDDCLK_posedge,
        TimingData     => Tmkr_LEDDADDR2_LEDDCLK_posedge,
        TestSignal     => LEDDADDR2_ipd,
        TestSignalName => "LEDDADDR2",
        TestDelay      => 0 ns,
        RefSignal      => LEDDCLK_ipd,
        RefSignalName  => "LEDDCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_LEDDADDR2_LEDDCLK_posedge_posedge,
        SetupLow       => tsetup_LEDDADDR2_LEDDCLK_negedge_posedge,
        HoldLow        => thold_LEDDADDR2_LEDDCLK_posedge_posedge,
        HoldHigh       => thold_LEDDADDR2_LEDDCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_LEDDA_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
		
		      VitalSetupHoldCheck (
        Violation      => Tviol_LEDDADDR3_LEDDCLK_posedge,
        TimingData     => Tmkr_LEDDADDR3_LEDDCLK_posedge,
        TestSignal     => LEDDADDR3_ipd,
        TestSignalName => "LEDDADDR3",
        TestDelay      => 0 ns,
        RefSignal      => LEDDCLK_ipd,
        RefSignalName  => "LEDDCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_LEDDADDR3_LEDDCLK_posedge_posedge,
        SetupLow       => tsetup_LEDDADDR3_LEDDCLK_negedge_posedge,
        HoldLow        => thold_LEDDADDR3_LEDDCLK_posedge_posedge,
        HoldHigh       => thold_LEDDADDR3_LEDDCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_LEDDA_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);		 
		
		   VitalSetupHoldCheck (
        Violation      => Tviol_LEDDDAT0_LEDDCLK_posedge,
        TimingData     => Tmkr_LEDDDAT0_LEDDCLK_posedge,
        TestSignal     => LEDDDAT0_ipd,
        TestSignalName => "LEDDDAT0",
        TestDelay      => 0 ns,
        RefSignal      => LEDDCLK_ipd,
        RefSignalName  => "LEDDCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_LEDDDAT0_LEDDCLK_posedge_posedge,
        SetupLow       => tsetup_LEDDDAT0_LEDDCLK_negedge_posedge,
        HoldLow        => thold_LEDDDAT0_LEDDCLK_posedge_posedge,
        HoldHigh       => thold_LEDDDAT0_LEDDCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_LEDDA_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
		
		   VitalSetupHoldCheck (
        Violation      => Tviol_LEDDDAT1_LEDDCLK_posedge,
        TimingData     => Tmkr_LEDDDAT1_LEDDCLK_posedge,
        TestSignal     => LEDDDAT1_ipd,
        TestSignalName => "LEDDDAT1",
        TestDelay      => 0 ns,
        RefSignal      => LEDDCLK_ipd,
        RefSignalName  => "LEDDCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_LEDDDAT1_LEDDCLK_posedge_posedge,
        SetupLow       => tsetup_LEDDDAT1_LEDDCLK_negedge_posedge,
        HoldLow        => thold_LEDDDAT1_LEDDCLK_posedge_posedge,
        HoldHigh       => thold_LEDDDAT1_LEDDCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_LEDDA_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
		
		   VitalSetupHoldCheck (
        Violation      => Tviol_LEDDDAT2_LEDDCLK_posedge,
        TimingData     => Tmkr_LEDDDAT2_LEDDCLK_posedge,
        TestSignal     => LEDDDAT2_ipd,
        TestSignalName => "LEDDDAT2",
        TestDelay      => 0 ns,
        RefSignal      => LEDDCLK_ipd,
        RefSignalName  => "LEDDCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_LEDDDAT2_LEDDCLK_posedge_posedge,
        SetupLow       => tsetup_LEDDDAT2_LEDDCLK_negedge_posedge,
        HoldLow        => thold_LEDDDAT2_LEDDCLK_posedge_posedge,
        HoldHigh       => thold_LEDDDAT2_LEDDCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_LEDDA_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
		
		
		   VitalSetupHoldCheck (
        Violation      => Tviol_LEDDDAT3_LEDDCLK_posedge,
        TimingData     => Tmkr_LEDDDAT3_LEDDCLK_posedge,
        TestSignal     => LEDDDAT3_ipd,
        TestSignalName => "LEDDDAT3",
        TestDelay      => 0 ns,
        RefSignal      => LEDDCLK_ipd,
        RefSignalName  => "LEDDCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_LEDDDAT3_LEDDCLK_posedge_posedge,
        SetupLow       => tsetup_LEDDDAT3_LEDDCLK_negedge_posedge,
        HoldLow        => thold_LEDDDAT3_LEDDCLK_posedge_posedge,
        HoldHigh       => thold_LEDDDAT3_LEDDCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_LEDDA_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
		
		
		   VitalSetupHoldCheck (
        Violation      => Tviol_LEDDDAT4_LEDDCLK_posedge,
        TimingData     => Tmkr_LEDDDAT4_LEDDCLK_posedge,
        TestSignal     => LEDDDAT4_ipd,
        TestSignalName => "LEDDDAT4",
        TestDelay      => 0 ns,
        RefSignal      => LEDDCLK_ipd,
        RefSignalName  => "LEDDCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_LEDDDAT4_LEDDCLK_posedge_posedge,
        SetupLow       => tsetup_LEDDDAT4_LEDDCLK_negedge_posedge,
        HoldLow        => thold_LEDDDAT4_LEDDCLK_posedge_posedge,
        HoldHigh       => thold_LEDDDAT4_LEDDCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_LEDDA_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
		
		
		   VitalSetupHoldCheck (
        Violation      => Tviol_LEDDDAT5_LEDDCLK_posedge,
        TimingData     => Tmkr_LEDDDAT5_LEDDCLK_posedge,
        TestSignal     => LEDDDAT5_ipd,
        TestSignalName => "LEDDDAT5",
        TestDelay      => 0 ns,
        RefSignal      => LEDDCLK_ipd,
        RefSignalName  => "LEDDCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_LEDDDAT5_LEDDCLK_posedge_posedge,
        SetupLow       => tsetup_LEDDDAT5_LEDDCLK_negedge_posedge,
        HoldLow        => thold_LEDDDAT5_LEDDCLK_posedge_posedge,
        HoldHigh       => thold_LEDDDAT5_LEDDCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_LEDDA_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
		
		
		   VitalSetupHoldCheck (
        Violation      => Tviol_LEDDDAT6_LEDDCLK_posedge,
        TimingData     => Tmkr_LEDDDAT6_LEDDCLK_posedge,
        TestSignal     => LEDDDAT6_ipd,
        TestSignalName => "LEDDDAT6",
        TestDelay      => 0 ns,
        RefSignal      => LEDDCLK_ipd,
        RefSignalName  => "LEDDCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_LEDDDAT6_LEDDCLK_posedge_posedge,
        SetupLow       => tsetup_LEDDDAT6_LEDDCLK_negedge_posedge,
        HoldLow        => thold_LEDDDAT6_LEDDCLK_posedge_posedge,
        HoldHigh       => thold_LEDDDAT6_LEDDCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_LEDDA_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
		
		
		   VitalSetupHoldCheck (
        Violation      => Tviol_LEDDDAT7_LEDDCLK_posedge,
        TimingData     => Tmkr_LEDDDAT7_LEDDCLK_posedge,
        TestSignal     => LEDDDAT7_ipd,
        TestSignalName => "LEDDDAT7",
        TestDelay      => 0 ns,
        RefSignal      => LEDDCLK_ipd,
        RefSignalName  => "LEDDCLK",
        RefDelay       => 0 ns,
        SetupHigh      => tsetup_LEDDDAT7_LEDDCLK_posedge_posedge,
        SetupLow       => tsetup_LEDDDAT7_LEDDCLK_negedge_posedge,
        HoldLow        => thold_LEDDDAT7_LEDDCLK_posedge_posedge,
        HoldHigh       => thold_LEDDDAT7_LEDDCLK_negedge_posedge,
        CheckEnabled   => true,
        RefTransition  => 'R',
        HeaderMsg      => "/SB_LEDDA_IP",
        Xon            => Xon,
        MsgOn          => MsgOn,
        MsgSeverity    => warning);	
end if; 		
----------------------
  --  Path Delay Section
  ----------------------
		
		    VitalPathDelay01 (
      OutSignal     => LEDDON,
      GlitchData    => LEDDON_GlitchData,
      OutSignalName => "LEDDON",
      OutTemp       => LEDDON_zd,
      Paths         => (0 => (LEDDCLK_ipd'last_event, tpd_LEDDCLK_LEDDON_posedge, true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);	
	    VitalPathDelay01 (
      OutSignal     => PWMOUT0,
      GlitchData    => PWMOUT0_GlitchData,
      OutSignalName => "PWMOUT0",
      OutTemp       => PWMOUT0_zd,
      Paths         => (0 => (LEDDCLK_ipd'last_event, tpd_LEDDCLK_PWMOUT0_posedge, true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);
	  
	     VitalPathDelay01 (
      OutSignal     => PWMOUT1,
      GlitchData    => PWMOUT1_GlitchData,
      OutSignalName => "PWMOUT1",
      OutTemp       => PWMOUT1_zd,
      Paths         => (0 => (LEDDCLK_ipd'last_event, tpd_LEDDCLK_PWMOUT1_posedge, true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);
	     VitalPathDelay01 (
      OutSignal     => PWMOUT2,
      GlitchData    => PWMOUT2_GlitchData,
      OutSignalName => "PWMOUT2",
      OutTemp       => PWMOUT2_zd,
      Paths         => (0 => (LEDDCLK_ipd'last_event, tpd_LEDDCLK_PWMOUT2_posedge, true)),
      Mode          => OnEvent,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning); 
	
end process VITALBehavior;
end 	SB_LEDDA_IP_V; 

--------------------------------------------
--------SMCCLK (20MHz Internal Clock) -----
-------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
library ieee;
use ieee.VITAL_Timing.all;
    
    
entity SMCCLK is
	Port (  CLK : out  std_logic ); 
end SMCCLK;

architecture SMCCLK_ARCH of SMCCLK is
	signal smc_clk :std_logic:='0';
begin

	process(smc_clk)
	begin 
		smc_clk<= not (smc_clk) after 25 ns;
	end process;

	CLK <= smc_clk;
 
end SMCCLK_ARCH; 

---------------------------------------------------
---- SB_SPRAM256KA --------------------------------
---------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
library ieee;
use ieee.VITAL_Timing.all; 

entity SB_SPRAM256KA is
	
		generic (	
		----------------------------------------------------------------------------------
		--VITAL PARAMETER
		---------------------------------------------------------------------------------
		TimingChecksOn  : boolean := true;
		Xon   		: boolean := true;
	        MsgOn 		: boolean := false;
		-- VITAL port delay
	        tipd_CLOCK  	: VitalDelayType01                   := ( 0 ns, 0 ns);
        	tipd_CHIPSELECT : VitalDelayType01                   := ( 0 ns, 0 ns);
		tipd_WREN    	: VitalDelayType01                   := ( 0 ns, 0 ns);
		tipd_STANDBY    : VitalDelayType01                   := ( 0 ns, 0 ns);
		tipd_SLEEP    	: VitalDelayType01                   := ( 0 ns, 0 ns);
		tipd_POWEROFF   : VitalDelayType01                   := ( 0 ns, 0 ns);
           	tipd_ADDRESS	: VitalDelayArrayType01(13 downto 0)  := (others => (0 ns, 0 ns));
           	tipd_DATAIN	: VitalDelayArrayType01(15 downto 0)  := (others => (0 ns, 0 ns));
           	tipd_MASKWREN	: VitalDelayArrayType01(3 downto 0)  := (others => (0 ns, 0 ns));
	         --- VITAL path delay
		--  VITAL clk-to-output path delay
		tpd_CLOCK_DATAOUT_posedge 		: VitalDelayArrayType01(15 downto 0) := (others => (0.000 ns, 0.000 ns));
       		tpd_SLEEP_DATAOUT_posedge 		: VitalDelayArrayType01(15 downto 0) :=(others => (0.000 ns, 0.000 ns));
		--- VITAL setup time
		tsetup_ADDRESS_CLOCK_negedge_posedge   	: VitalDelayArrayType(13 downto 0) := (others => 0 ns );
	        tsetup_ADDRESS_CLOCK_posedge_posedge   	: VitalDelayArrayType(13 downto 0) := (others => 0 ns );
	        tsetup_DATAIN_CLOCK_negedge_posedge    	: VitalDelayArrayType(15 downto 0) := (others => 0 ns );
	        tsetup_DATAIN_CLOCK_posedge_posedge    	: VitalDelayArrayType(15 downto 0) := (others => 0 ns );
		tsetup_MASKWREN_CLOCK_negedge_posedge  	: VitalDelayArrayType(3 downto 0) := (others => 0 ns );
	        tsetup_MASKWREN_CLOCK_posedge_posedge  	: VitalDelayArrayType(3 downto 0) := (others => 0 ns );

       		tsetup_WREN_CLOCK_negedge_posedge 	: VitalDelayType := 0 ns;
	        tsetup_WREN_CLOCK_posedge_posedge 	: VitalDelayType := 0 ns;
	        tsetup_CHIPSELECT_CLOCK_posedge_posedge	: VitalDelayType := 0 ns;
	        tsetup_CHIPSELECT_CLOCK_negedge_posedge	: VitalDelayType := 0 ns;

		tsetup_STANDBY_CLOCK_negedge_posedge   	: VitalDelayType := 0 ns;
           	tsetup_STANDBY_CLOCK_posedge_posedge   	: VitalDelayType := 0 ns;
		tsetup_SLEEP_CLOCK_negedge_posedge 	: VitalDelayType := 0 ns;
           	tsetup_SLEEP_CLOCK_posedge_posedge 	: VitalDelayType := 0 ns;

		--- VITAL hold time
		thold_ADDRESS_CLOCK_negedge_posedge   	: VitalDelayArrayType(13 downto 0) := (others => 0 ns );
	        thold_ADDRESS_CLOCK_posedge_posedge   	: VitalDelayArrayType(13 downto 0) := (others => 0 ns );
	        thold_DATAIN_CLOCK_negedge_posedge    	: VitalDelayArrayType(15 downto 0) := (others => 0 ns );
	        thold_DATAIN_CLOCK_posedge_posedge    	: VitalDelayArrayType(15 downto 0) := (others => 0 ns );
		thold_MASKWREN_CLOCK_negedge_posedge  	: VitalDelayArrayType(3 downto 0) := (others => 0 ns );
	        thold_MASKWREN_CLOCK_posedge_posedge  	: VitalDelayArrayType(3 downto 0) := (others => 0 ns );

       		thold_WREN_CLOCK_negedge_posedge 	: VitalDelayType := 0 ns;
	        thold_WREN_CLOCK_posedge_posedge 	: VitalDelayType := 0 ns;
	        thold_CHIPSELECT_CLOCK_posedge_posedge	: VitalDelayType := 0 ns;
	        thold_CHIPSELECT_CLOCK_negedge_posedge	: VitalDelayType := 0 ns;

		thold_STANDBY_CLOCK_negedge_posedge   	: VitalDelayType := 0 ns;
           	thold_STANDBY_CLOCK_posedge_posedge   	: VitalDelayType := 0 ns;
		thold_SLEEP_CLOCK_negedge_posedge 	: VitalDelayType := 0 ns;
		thold_SLEEP_CLOCK_posedge_posedge 	: VitalDelayType := 0 ns
		);


	Port (  CLOCK 	: in std_logic ;	
		ADDRESS : in std_logic_vector(13 downto 0); 
		DATAIN  : in std_logic_vector(15 downto 0); 
		MASKWREN : in std_logic_vector(3 downto 0); 
		WREN	: in std_logic; 
		CHIPSELECT: in std_logic ; 
		STANDBY	: in std_logic := 'L' ; 
		SLEEP	: in std_logic := 'L' ; 
		POWEROFF: in std_logic := 'H' ;		--  Note : 1'b0 to POWEROFF RAM  , 1'b1 to POWERON RAM block at wrapper level.  
		DATAOUT	: out std_logic_vector(15 downto 0)		
	     ); 

	attribute VITAL_LEVEL0 of  SB_SPRAM256KA : entity is true;	

end SB_SPRAM256KA;


architecture SB_SPRAM256KA_V of SB_SPRAM256KA is

attribute VITAL_LEVEL0 of
    SB_SPRAM256KA_V : architecture is true;


component sadslspk4s1p16384x16m16b4w1c0p1d0t0 is
	port (
		CLK 	: in std_logic ;	
		ADR 	: in std_logic_vector(13 downto 0); 
		D  	: in std_logic_vector(15 downto 0); 
		WEM 	: in std_logic_vector(15 downto 0); 
		WE	: in std_logic; 
		ME	: in std_logic ; 
		LS	: in std_logic; 
		DS	: in std_logic; 
		SD	: in std_logic; 
		Q	: out std_logic_vector(15 downto 0);
		TEST1	: in  std_logic ;
		RME	: in  std_logic; 
		RM	: in   std_logic_vector(3 downto 0)
		);
end component;

	--- VITAL Signals   
	signal ADDRESS_ipd : std_logic_vector(13 downto 0)  := (others => 'X');   
	signal DATAIN_ipd : std_logic_vector(15 downto 0)  := (others => 'X');   
	signal MASKWREN_ipd : std_logic_vector(3 downto 0)  := (others => 'X');   
	signal CLOCK_ipd  : std_logic                    := 'X';
	signal WREN_ipd : std_logic                    := 'X';
	signal CHIPSELECT_ipd    : std_logic                    := 'X';
	signal STANDBY_ipd  : std_logic                    := 'X';  
	signal SLEEP_ipd  : std_logic                    := 'X';  
	signal POWEROFF_ipd  : std_logic                    := 'X';  
	signal not_poweroff  : std_logic :='X'; 

	signal DATAOUT_zd : std_logic_vector(15 downto 0)  := (others => 'X');   

 	-- Functional Signals. 

	signal maskwem	: std_logic_vector(15 downto 0) := (others => 'X');  


begin 	

	---------------------
	--  Input Wire Delay
	---------------------
	WireDelay : block
	begin
	  ADDRESS_DELAY : for i in 13 downto 0 generate
	     VitalWireDelay (ADDRESS_ipd(i), ADDRESS(i), tipd_ADDRESS(i));
	  end generate ADDRESS_DELAY;
  	  DATAIN_DELAY : for i in 15 downto 0 generate
	     VitalWireDelay (DATAIN_ipd(i), DATAIN(i), tipd_DATAIN(i));
	  end generate DATAIN_DELAY;
  	  MASKWREN_DELAY : for i in 3 downto 0 generate
	     VitalWireDelay (MASKWREN_ipd(i), MASKWREN(i), tipd_MASKWREN(i));
	  end generate MASKWREN_DELAY;
	  VitalWireDelay (CLOCK_ipd, CLOCK, tipd_CLOCK);
	  VitalWireDelay (WREN_ipd, WREN, tipd_WREN);
	  VitalWireDelay (CHIPSELECT_ipd, CHIPSELECT, tipd_CHIPSELECT);
	  VitalWireDelay (STANDBY_ipd, STANDBY, tipd_STANDBY);
	  VitalWireDelay (SLEEP_ipd, SLEEP, tipd_SLEEP);
	  VitalWireDelay (POWEROFF_ipd, POWEROFF, tipd_POWEROFF);

	end block WireDelay;
	
	VITALBehavior : block
	begin
	---------------------
	--  Timing Checks
	---------------------
	TimingChecks : process (ADDRESS_ipd, DATAIN_ipd, MASKWREN_ipd, CLOCK_ipd, WREN_ipd, CHIPSELECT_ipd, STANDBY_ipd, SLEEP_ipd, POWEROFF_ipd)

	variable Tviol_ADDRESS_CLOCK_posedge : std_logic_vector(13 downto 0) :=(others => '0');
	variable Tviol_DATAIN_CLOCK_posedge : std_logic_vector(15 downto 0) :=(others => '0');
	variable Tviol_MASKWREN_CLOCK_posedge : std_logic_vector(3 downto 0) :=(others => '0');
	variable Tviol_WREN_CLOCK_posedge  : std_logic := '0';
	variable Tviol_CHIPSELECT_CLOCK_posedge  : std_logic := '0';
	variable Tviol_STANDBY_CLOCK_posedge  : std_logic := '0';
	variable Tviol_SLEEP_CLOCK_posedge  : std_logic := '0';


	variable Tmkr_ADDRESS0_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_ADDRESS1_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_ADDRESS2_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_ADDRESS3_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_ADDRESS4_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_ADDRESS5_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_ADDRESS6_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_ADDRESS7_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_ADDRESS8_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_ADDRESS9_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_ADDRESS10_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_ADDRESS11_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_ADDRESS12_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_ADDRESS13_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;

	variable Tmkr_DATAIN0_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DATAIN1_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DATAIN2_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DATAIN3_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DATAIN4_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DATAIN5_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DATAIN6_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DATAIN7_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DATAIN8_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DATAIN9_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DATAIN10_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DATAIN11_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DATAIN12_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DATAIN13_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DATAIN14_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DATAIN15_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;

	variable Tmkr_MASKWREN0_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MASKWREN1_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MASKWREN2_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MASKWREN3_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;

	variable Tmkr_WREN_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_CHIPSELECT_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_SLEEP_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_STANDBY_CLOCK_posedge : VitalTimingDataType := VitalTimingDataInit;

	variable PViol_CLOCK : std_logic := '0'; 
	variable PInfo_CLOCK : VitalPeriodDataType;

	variable Violation     : std_logic  := '0';

	begin

	    if (TimingChecksOn) then
	      VitalSetupHoldCheck (
		Violation      => Tviol_ADDRESS_CLOCK_posedge(0),
		TimingData     => Tmkr_ADDRESS0_CLOCK_posedge,
		TestSignal     => ADDRESS_ipd(0),
		TestSignalName => "ADDRESS(0)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_ADDRESS_CLOCK_posedge_posedge(0),
		SetupLow       => tsetup_ADDRESS_CLOCK_negedge_posedge(0),
		HoldLow        => thold_ADDRESS_CLOCK_posedge_posedge(0),
		HoldHigh       => thold_ADDRESS_CLOCK_negedge_posedge(0),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_ADDRESS_CLOCK_posedge(1),
		TimingData     => Tmkr_ADDRESS1_CLOCK_posedge,
		TestSignal     => ADDRESS_ipd(1),
		TestSignalName => "ADDRESS(1)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_ADDRESS_CLOCK_posedge_posedge(1),
		SetupLow       => tsetup_ADDRESS_CLOCK_negedge_posedge(1),
		HoldLow        => thold_ADDRESS_CLOCK_posedge_posedge(1),
		HoldHigh       => thold_ADDRESS_CLOCK_negedge_posedge(1),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
			      VitalSetupHoldCheck (
		Violation      => Tviol_ADDRESS_CLOCK_posedge(2),
		TimingData     => Tmkr_ADDRESS2_CLOCK_posedge,
		TestSignal     => ADDRESS_ipd(2),
		TestSignalName => "ADDRESS(2)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_ADDRESS_CLOCK_posedge_posedge(2),
		SetupLow       => tsetup_ADDRESS_CLOCK_negedge_posedge(2),
		HoldLow        => thold_ADDRESS_CLOCK_posedge_posedge(2),
		HoldHigh       => thold_ADDRESS_CLOCK_negedge_posedge(2),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_ADDRESS_CLOCK_posedge(3),
		TimingData     => Tmkr_ADDRESS3_CLOCK_posedge,
		TestSignal     => ADDRESS_ipd(3),
		TestSignalName => "ADDRESS(3)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_ADDRESS_CLOCK_posedge_posedge(3),
		SetupLow       => tsetup_ADDRESS_CLOCK_negedge_posedge(3),
		HoldLow        => thold_ADDRESS_CLOCK_posedge_posedge(3),
		HoldHigh       => thold_ADDRESS_CLOCK_negedge_posedge(3),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	     VitalSetupHoldCheck (
		Violation      => Tviol_ADDRESS_CLOCK_posedge(4),
		TimingData     => Tmkr_ADDRESS4_CLOCK_posedge,
		TestSignal     => ADDRESS_ipd(4),
		TestSignalName => "ADDRESS(4)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_ADDRESS_CLOCK_posedge_posedge(4),
		SetupLow       => tsetup_ADDRESS_CLOCK_negedge_posedge(4),
		HoldLow        => thold_ADDRESS_CLOCK_posedge_posedge(4),
		HoldHigh       => thold_ADDRESS_CLOCK_negedge_posedge(4),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_ADDRESS_CLOCK_posedge(5),
		TimingData     => Tmkr_ADDRESS5_CLOCK_posedge,
		TestSignal     => ADDRESS_ipd(5),
		TestSignalName => "ADDRESS(5)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_ADDRESS_CLOCK_posedge_posedge(5),
		SetupLow       => tsetup_ADDRESS_CLOCK_negedge_posedge(5),
		HoldLow        => thold_ADDRESS_CLOCK_posedge_posedge(5),
		HoldHigh       => thold_ADDRESS_CLOCK_negedge_posedge(5),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_ADDRESS_CLOCK_posedge(6),
		TimingData     => Tmkr_ADDRESS6_CLOCK_posedge,
		TestSignal     => ADDRESS_ipd(6),
		TestSignalName => "ADDRESS(6)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_ADDRESS_CLOCK_posedge_posedge(6),
		SetupLow       => tsetup_ADDRESS_CLOCK_negedge_posedge(6),
		HoldLow        => thold_ADDRESS_CLOCK_posedge_posedge(6),
		HoldHigh       => thold_ADDRESS_CLOCK_negedge_posedge(6),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_ADDRESS_CLOCK_posedge(7),
		TimingData     => Tmkr_ADDRESS7_CLOCK_posedge,
		TestSignal     => ADDRESS_ipd(7),
		TestSignalName => "ADDRESS(7)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_ADDRESS_CLOCK_posedge_posedge(7),
		SetupLow       => tsetup_ADDRESS_CLOCK_negedge_posedge(7),
		HoldLow        => thold_ADDRESS_CLOCK_posedge_posedge(7),
		HoldHigh       => thold_ADDRESS_CLOCK_negedge_posedge(7),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_ADDRESS_CLOCK_posedge(8),
		TimingData     => Tmkr_ADDRESS8_CLOCK_posedge,
		TestSignal     => ADDRESS_ipd(8),
		TestSignalName => "ADDRESS(8)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_ADDRESS_CLOCK_posedge_posedge(8),
		SetupLow       => tsetup_ADDRESS_CLOCK_negedge_posedge(8),
		HoldLow        => thold_ADDRESS_CLOCK_posedge_posedge(8),
		HoldHigh       => thold_ADDRESS_CLOCK_negedge_posedge(8),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_ADDRESS_CLOCK_posedge(9),
		TimingData     => Tmkr_ADDRESS9_CLOCK_posedge,
		TestSignal     => ADDRESS_ipd(9),
		TestSignalName => "ADDRESS(9)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_ADDRESS_CLOCK_posedge_posedge(9),
		SetupLow       => tsetup_ADDRESS_CLOCK_negedge_posedge(9),
		HoldLow        => thold_ADDRESS_CLOCK_posedge_posedge(9),
		HoldHigh       => thold_ADDRESS_CLOCK_negedge_posedge(9),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_ADDRESS_CLOCK_posedge(10),
		TimingData     => Tmkr_ADDRESS10_CLOCK_posedge,
		TestSignal     => ADDRESS_ipd(10),
		TestSignalName => "ADDRESS(10)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_ADDRESS_CLOCK_posedge_posedge(10),
		SetupLow       => tsetup_ADDRESS_CLOCK_negedge_posedge(10),
		HoldLow        => thold_ADDRESS_CLOCK_posedge_posedge(10),
		HoldHigh       => thold_ADDRESS_CLOCK_negedge_posedge(10),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_ADDRESS_CLOCK_posedge(11),
		TimingData     => Tmkr_ADDRESS11_CLOCK_posedge,
		TestSignal     => ADDRESS_ipd(11),
		TestSignalName => "ADDRESS(11)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_ADDRESS_CLOCK_posedge_posedge(11),
		SetupLow       => tsetup_ADDRESS_CLOCK_negedge_posedge(11),
		HoldLow        => thold_ADDRESS_CLOCK_posedge_posedge(11),
		HoldHigh       => thold_ADDRESS_CLOCK_negedge_posedge(11),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_ADDRESS_CLOCK_posedge(12),
		TimingData     => Tmkr_ADDRESS12_CLOCK_posedge,
		TestSignal     => ADDRESS_ipd(12),
		TestSignalName => "ADDRESS(12)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_ADDRESS_CLOCK_posedge_posedge(12),
		SetupLow       => tsetup_ADDRESS_CLOCK_negedge_posedge(12),
		HoldLow        => thold_ADDRESS_CLOCK_posedge_posedge(12),
		HoldHigh       => thold_ADDRESS_CLOCK_negedge_posedge(12),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_ADDRESS_CLOCK_posedge(13),
		TimingData     => Tmkr_ADDRESS13_CLOCK_posedge,
		TestSignal     => ADDRESS_ipd(13),
		TestSignalName => "ADDRESS(13)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_ADDRESS_CLOCK_posedge_posedge(13),
		SetupLow       => tsetup_ADDRESS_CLOCK_negedge_posedge(13),
		HoldLow        => thold_ADDRESS_CLOCK_posedge_posedge(13),
		HoldHigh       => thold_ADDRESS_CLOCK_negedge_posedge(13),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	-- DATAIN
	    VitalSetupHoldCheck (
		Violation      => Tviol_DATAIN_CLOCK_posedge(0),
		TimingData     => Tmkr_DATAIN0_CLOCK_posedge,
		TestSignal     => DATAIN_ipd(0),
		TestSignalName => "DATAIN(0)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_DATAIN_CLOCK_posedge_posedge(0),
		SetupLow       => tsetup_DATAIN_CLOCK_negedge_posedge(0),
		HoldLow        => thold_DATAIN_CLOCK_posedge_posedge(0),
		HoldHigh       => thold_DATAIN_CLOCK_negedge_posedge(0),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_DATAIN_CLOCK_posedge(1),
		TimingData     => Tmkr_DATAIN1_CLOCK_posedge,
		TestSignal     => DATAIN_ipd(1),
		TestSignalName => "DATAIN(1)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_DATAIN_CLOCK_posedge_posedge(1),
		SetupLow       => tsetup_DATAIN_CLOCK_negedge_posedge(1),
		HoldLow        => thold_DATAIN_CLOCK_posedge_posedge(1),
		HoldHigh       => thold_DATAIN_CLOCK_negedge_posedge(1),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
			      VitalSetupHoldCheck (
		Violation      => Tviol_DATAIN_CLOCK_posedge(2),
		TimingData     => Tmkr_DATAIN2_CLOCK_posedge,
		TestSignal     => DATAIN_ipd(2),
		TestSignalName => "DATAIN(2)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_DATAIN_CLOCK_posedge_posedge(2),
		SetupLow       => tsetup_DATAIN_CLOCK_negedge_posedge(2),
		HoldLow        => thold_DATAIN_CLOCK_posedge_posedge(2),
		HoldHigh       => thold_DATAIN_CLOCK_negedge_posedge(2),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_DATAIN_CLOCK_posedge(3),
		TimingData     => Tmkr_DATAIN3_CLOCK_posedge,
		TestSignal     => DATAIN_ipd(3),
		TestSignalName => "DATAIN(3)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_DATAIN_CLOCK_posedge_posedge(3),
		SetupLow       => tsetup_DATAIN_CLOCK_negedge_posedge(3),
		HoldLow        => thold_DATAIN_CLOCK_posedge_posedge(3),
		HoldHigh       => thold_DATAIN_CLOCK_negedge_posedge(3),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	     VitalSetupHoldCheck (
		Violation      => Tviol_DATAIN_CLOCK_posedge(4),
		TimingData     => Tmkr_DATAIN4_CLOCK_posedge,
		TestSignal     => DATAIN_ipd(4),
		TestSignalName => "DATAIN(4)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_DATAIN_CLOCK_posedge_posedge(4),
		SetupLow       => tsetup_DATAIN_CLOCK_negedge_posedge(4),
		HoldLow        => thold_DATAIN_CLOCK_posedge_posedge(4),
		HoldHigh       => thold_DATAIN_CLOCK_negedge_posedge(4),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_DATAIN_CLOCK_posedge(5),
		TimingData     => Tmkr_DATAIN5_CLOCK_posedge,
		TestSignal     => DATAIN_ipd(5),
		TestSignalName => "DATAIN(5)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_DATAIN_CLOCK_posedge_posedge(5),
		SetupLow       => tsetup_DATAIN_CLOCK_negedge_posedge(5),
		HoldLow        => thold_DATAIN_CLOCK_posedge_posedge(5),
		HoldHigh       => thold_DATAIN_CLOCK_negedge_posedge(5),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_DATAIN_CLOCK_posedge(6),
		TimingData     => Tmkr_DATAIN6_CLOCK_posedge,
		TestSignal     => DATAIN_ipd(6),
		TestSignalName => "DATAIN(6)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_DATAIN_CLOCK_posedge_posedge(6),
		SetupLow       => tsetup_DATAIN_CLOCK_negedge_posedge(6),
		HoldLow        => thold_DATAIN_CLOCK_posedge_posedge(6),
		HoldHigh       => thold_DATAIN_CLOCK_negedge_posedge(6),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_DATAIN_CLOCK_posedge(7),
		TimingData     => Tmkr_DATAIN7_CLOCK_posedge,
		TestSignal     => DATAIN_ipd(7),
		TestSignalName => "DATAIN(7)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_DATAIN_CLOCK_posedge_posedge(7),
		SetupLow       => tsetup_DATAIN_CLOCK_negedge_posedge(7),
		HoldLow        => thold_DATAIN_CLOCK_posedge_posedge(7),
		HoldHigh       => thold_DATAIN_CLOCK_negedge_posedge(7),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_DATAIN_CLOCK_posedge(8),
		TimingData     => Tmkr_DATAIN8_CLOCK_posedge,
		TestSignal     => DATAIN_ipd(8),
		TestSignalName => "DATAIN(8)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_DATAIN_CLOCK_posedge_posedge(8),
		SetupLow       => tsetup_DATAIN_CLOCK_negedge_posedge(8),
		HoldLow        => thold_DATAIN_CLOCK_posedge_posedge(8),
		HoldHigh       => thold_DATAIN_CLOCK_negedge_posedge(8),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_DATAIN_CLOCK_posedge(9),
		TimingData     => Tmkr_DATAIN9_CLOCK_posedge,
		TestSignal     => DATAIN_ipd(9),
		TestSignalName => "DATAIN(9)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_DATAIN_CLOCK_posedge_posedge(9),
		SetupLow       => tsetup_DATAIN_CLOCK_negedge_posedge(9),
		HoldLow        => thold_DATAIN_CLOCK_posedge_posedge(9),
		HoldHigh       => thold_DATAIN_CLOCK_negedge_posedge(9),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_DATAIN_CLOCK_posedge(10),
		TimingData     => Tmkr_DATAIN10_CLOCK_posedge,
		TestSignal     => DATAIN_ipd(10),
		TestSignalName => "DATAIN(10)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_DATAIN_CLOCK_posedge_posedge(10),
		SetupLow       => tsetup_DATAIN_CLOCK_negedge_posedge(10),
		HoldLow        => thold_DATAIN_CLOCK_posedge_posedge(10),
		HoldHigh       => thold_DATAIN_CLOCK_negedge_posedge(10),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_DATAIN_CLOCK_posedge(11),
		TimingData     => Tmkr_DATAIN11_CLOCK_posedge,
		TestSignal     => DATAIN_ipd(11),
		TestSignalName => "DATAIN(11)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_DATAIN_CLOCK_posedge_posedge(11),
		SetupLow       => tsetup_DATAIN_CLOCK_negedge_posedge(11),
		HoldLow        => thold_DATAIN_CLOCK_posedge_posedge(11),
		HoldHigh       => thold_DATAIN_CLOCK_negedge_posedge(11),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	     VitalSetupHoldCheck (
		Violation      => Tviol_DATAIN_CLOCK_posedge(12),
		TimingData     => Tmkr_DATAIN12_CLOCK_posedge,
		TestSignal     => DATAIN_ipd(12),
		TestSignalName => "DATAIN(12)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_DATAIN_CLOCK_posedge_posedge(12),
		SetupLow       => tsetup_DATAIN_CLOCK_negedge_posedge(12),
		HoldLow        => thold_DATAIN_CLOCK_posedge_posedge(12),
		HoldHigh       => thold_DATAIN_CLOCK_negedge_posedge(12),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_DATAIN_CLOCK_posedge(13),
		TimingData     => Tmkr_DATAIN13_CLOCK_posedge,
		TestSignal     => DATAIN_ipd(13),
		TestSignalName => "DATAIN(13)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_DATAIN_CLOCK_posedge_posedge(13),
		SetupLow       => tsetup_DATAIN_CLOCK_negedge_posedge(13),
		HoldLow        => thold_DATAIN_CLOCK_posedge_posedge(13),
		HoldHigh       => thold_DATAIN_CLOCK_negedge_posedge(13),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	     VitalSetupHoldCheck (
		Violation      => Tviol_DATAIN_CLOCK_posedge(14),
		TimingData     => Tmkr_DATAIN14_CLOCK_posedge,
		TestSignal     => DATAIN_ipd(14),
		TestSignalName => "DATAIN(14)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_DATAIN_CLOCK_posedge_posedge(14),
		SetupLow       => tsetup_DATAIN_CLOCK_negedge_posedge(14),
		HoldLow        => thold_DATAIN_CLOCK_posedge_posedge(14),
		HoldHigh       => thold_DATAIN_CLOCK_negedge_posedge(14),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_DATAIN_CLOCK_posedge(15),
		TimingData     => Tmkr_DATAIN15_CLOCK_posedge,
		TestSignal     => DATAIN_ipd(15),
		TestSignalName => "DATAIN(15)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_DATAIN_CLOCK_posedge_posedge(15),
		SetupLow       => tsetup_DATAIN_CLOCK_negedge_posedge(15),
		HoldLow        => thold_DATAIN_CLOCK_posedge_posedge(15),
		HoldHigh       => thold_DATAIN_CLOCK_negedge_posedge(15),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	-- MASKWREN
	    VitalSetupHoldCheck (
		Violation      => Tviol_MASKWREN_CLOCK_posedge(0),
		TimingData     => Tmkr_MASKWREN0_CLOCK_posedge,
		TestSignal     => MASKWREN_ipd(0),
		TestSignalName => "MASKWREN(0)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASKWREN_CLOCK_posedge_posedge(0),
		SetupLow       => tsetup_MASKWREN_CLOCK_negedge_posedge(0),
		HoldLow        => thold_MASKWREN_CLOCK_posedge_posedge(0),
		HoldHigh       => thold_MASKWREN_CLOCK_negedge_posedge(0),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_MASKWREN_CLOCK_posedge(1),
		TimingData     => Tmkr_MASKWREN1_CLOCK_posedge,
		TestSignal     => MASKWREN_ipd(1),
		TestSignalName => "MASKWREN(1)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASKWREN_CLOCK_posedge_posedge(1),
		SetupLow       => tsetup_MASKWREN_CLOCK_negedge_posedge(1),
		HoldLow        => thold_MASKWREN_CLOCK_posedge_posedge(1),
		HoldHigh       => thold_MASKWREN_CLOCK_negedge_posedge(1),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	     VitalSetupHoldCheck (
		Violation      => Tviol_MASKWREN_CLOCK_posedge(2),
		TimingData     => Tmkr_MASKWREN2_CLOCK_posedge,
		TestSignal     => MASKWREN_ipd(2),
		TestSignalName => "MASKWREN(2)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASKWREN_CLOCK_posedge_posedge(2),
		SetupLow       => tsetup_MASKWREN_CLOCK_negedge_posedge(2),
		HoldLow        => thold_MASKWREN_CLOCK_posedge_posedge(2),
		HoldHigh       => thold_MASKWREN_CLOCK_negedge_posedge(2),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_MASKWREN_CLOCK_posedge(3),
		TimingData     => Tmkr_MASKWREN3_CLOCK_posedge,
		TestSignal     => MASKWREN_ipd(3),
		TestSignalName => "MASKWREN(3)",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_MASKWREN_CLOCK_posedge_posedge(3),
		SetupLow       => tsetup_MASKWREN_CLOCK_negedge_posedge(3),
		HoldLow        => thold_MASKWREN_CLOCK_posedge_posedge(3),
		HoldHigh       => thold_MASKWREN_CLOCK_negedge_posedge(3),
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	-- WREN

	      VitalSetupHoldCheck (
		Violation      => Tviol_WREN_CLOCK_posedge,
		TimingData     => Tmkr_WREN_CLOCK_posedge,
		TestSignal     => WREN_ipd,
		TestSignalName => "WREN",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_WREN_CLOCK_posedge_posedge,
		SetupLow       => tsetup_WREN_CLOCK_negedge_posedge,
		HoldLow        => thold_WREN_CLOCK_posedge_posedge,
		HoldHigh       => thold_WREN_CLOCK_negedge_posedge,
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_RAM40_4K",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		
	      VitalSetupHoldCheck (
		Violation      => Tviol_CHIPSELECT_CLOCK_posedge,
		TimingData     => Tmkr_CHIPSELECT_CLOCK_posedge,
		TestSignal     => CHIPSELECT_ipd,
		TestSignalName => "CHIPSELECT",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_CHIPSELECT_CLOCK_posedge_posedge,
		SetupLow       => tsetup_CHIPSELECT_CLOCK_negedge_posedge,
		HoldLow        => thold_CHIPSELECT_CLOCK_posedge_posedge,
		HoldHigh       => thold_CHIPSELECT_CLOCK_negedge_posedge,
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);
		       

	      VitalSetupHoldCheck (
		Violation      => Tviol_STANDBY_CLOCK_posedge,
		TimingData     => Tmkr_STANDBY_CLOCK_posedge,
		TestSignal     => STANDBY_ipd,
		TestSignalName => "STANDBY",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_STANDBY_CLOCK_posedge_posedge,
		SetupLow       => tsetup_STANDBY_CLOCK_negedge_posedge,
		HoldLow        => thold_STANDBY_CLOCK_posedge_posedge,
		HoldHigh       => thold_STANDBY_CLOCK_negedge_posedge,
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	      VitalSetupHoldCheck (
		Violation      => Tviol_SLEEP_CLOCK_posedge,
		TimingData     => Tmkr_SLEEP_CLOCK_posedge,
		TestSignal     => SLEEP_ipd,
		TestSignalName => "SLEEP",
		TestDelay      => 0 ns,
		RefSignal      => CLOCK_ipd,
		RefSignalName  => "CLOCK",
		RefDelay       => 0 ns,
		SetupHigh      => tsetup_SLEEP_CLOCK_posedge_posedge,
		SetupLow       => tsetup_SLEEP_CLOCK_negedge_posedge,
		HoldLow        => thold_SLEEP_CLOCK_posedge_posedge,
		HoldHigh       => thold_SLEEP_CLOCK_negedge_posedge,
		CheckEnabled   => true,
		RefTransition  => 'R',
		HeaderMsg      => "/SB_SPRAM256KA",
		Xon            => Xon,
		MsgOn          => MsgOn,
		MsgSeverity    => warning);

	    Violation  := Tviol_ADDRESS_CLOCK_posedge(0) or
			  Tviol_ADDRESS_CLOCK_posedge(1) or
			  Tviol_ADDRESS_CLOCK_posedge(2) or
	  		  Tviol_ADDRESS_CLOCK_posedge(3) or
	  		  Tviol_ADDRESS_CLOCK_posedge(4) or
	  		  Tviol_ADDRESS_CLOCK_posedge(5) or
	  		  Tviol_ADDRESS_CLOCK_posedge(6) or
			  Tviol_ADDRESS_CLOCK_posedge(7) or
			  Tviol_ADDRESS_CLOCK_posedge(8) or			  
			  Tviol_ADDRESS_CLOCK_posedge(9) or			  
			  Tviol_ADDRESS_CLOCK_posedge(10) or			  
	  		  Tviol_ADDRESS_CLOCK_posedge(11) or
			  Tviol_ADDRESS_CLOCK_posedge(12) or			  
			  Tviol_ADDRESS_CLOCK_posedge(13) or
			  Tviol_DATAIN_CLOCK_posedge(0) or	
  			  Tviol_DATAIN_CLOCK_posedge(1) or
			  Tviol_DATAIN_CLOCK_posedge(2) or
	  		  Tviol_DATAIN_CLOCK_posedge(3) or
	  		  Tviol_DATAIN_CLOCK_posedge(4) or
	  		  Tviol_DATAIN_CLOCK_posedge(5) or
	  		  Tviol_DATAIN_CLOCK_posedge(6) or
			  Tviol_DATAIN_CLOCK_posedge(7) or
			  Tviol_DATAIN_CLOCK_posedge(8) or			  
			  Tviol_DATAIN_CLOCK_posedge(9) or			  
			  Tviol_DATAIN_CLOCK_posedge(10) or			  
	  		  Tviol_DATAIN_CLOCK_posedge(11) or
			  Tviol_DATAIN_CLOCK_posedge(12) or			  
			  Tviol_DATAIN_CLOCK_posedge(13) or
			  Tviol_DATAIN_CLOCK_posedge(14) or
  			  Tviol_DATAIN_CLOCK_posedge(15) or
			  Tviol_MASKWREN_CLOCK_posedge(0) or	
  			  Tviol_MASKWREN_CLOCK_posedge(1) or
			  Tviol_MASKWREN_CLOCK_posedge(2) or
	  		  Tviol_MASKWREN_CLOCK_posedge(3) or
			  Tviol_WREN_CLOCK_posedge or
			  Tviol_CHIPSELECT_CLOCK_posedge or
			  Tviol_STANDBY_CLOCK_posedge or
			  Tviol_SLEEP_CLOCK_posedge ; 

		assert violation = '0'
			report " Incorrect due to Timing Violations\n"
		severity warning;

	    end if ;
    end process TimingChecks;

	----------------------------
	--- Behavioural section
	------------------------------

	maskwem <= ( MASKWREN_ipd(3) & MASKWREN_ipd(3) & MASKWREN_ipd(3) & MASKWREN_ipd(3) & MASKWREN_ipd(2) & MASKWREN_ipd(2) & MASKWREN(2) & MASKWREN_ipd(2) & MASKWREN_ipd(1) & MASKWREN_ipd(1) & MASKWREN_ipd(1) & MASKWREN_ipd(1) & MASKWREN_ipd(0) & MASKWREN_ipd(0) & MASKWREN_ipd(0) & MASKWREN_ipd(0) );

	not_poweroff <= not(POWEROFF_ipd); 

spram256k_core_inst :  sadslspk4s1p16384x16m16b4w1c0p1d0t0
	port map    	(
	        CLK => CLOCK_ipd, 
		ADR => ADDRESS_ipd, 
		D  	=> DATAIN_ipd, 
		WEM => maskwem, 
		WE	=> WREN_ipd, 
		ME	=> CHIPSELECT_ipd, 
		LS	=> STANDBY_ipd, 
		DS	=> SLEEP_ipd, 
		SD	=> not_poweroff, 
		Q	=> DATAOUT_zd, 
		TEST1 	=> '0', 
		RME	=> '0',
		RM	=> "0000"
		);

	------------------------- 
	--- Path delay section 
   	------------------------ 
	PathDelay : process(DATAOUT_zd)

	variable DATAOUT_GlitchData0  : VitalGlitchDataType;
	variable DATAOUT_GlitchData1  : VitalGlitchDataType;
	variable DATAOUT_GlitchData2  : VitalGlitchDataType;
	variable DATAOUT_GlitchData3  : VitalGlitchDataType;
	variable DATAOUT_GlitchData4  : VitalGlitchDataType;
	variable DATAOUT_GlitchData5  : VitalGlitchDataType;
	variable DATAOUT_GlitchData6  : VitalGlitchDataType;
	variable DATAOUT_GlitchData7  : VitalGlitchDataType;
	variable DATAOUT_GlitchData8  : VitalGlitchDataType;
	variable DATAOUT_GlitchData9  : VitalGlitchDataType;
	variable DATAOUT_GlitchData10 : VitalGlitchDataType;
	variable DATAOUT_GlitchData11 : VitalGlitchDataType;
	variable DATAOUT_GlitchData12 : VitalGlitchDataType;
	variable DATAOUT_GlitchData13 : VitalGlitchDataType;
	variable DATAOUT_GlitchData14 : VitalGlitchDataType;
	variable DATAOUT_GlitchData15 : VitalGlitchDataType;
	begin
	    VitalPathDelay01 (
	      OutSignal     => DATAOUT(0),
	      GlitchData    => DATAOUT_GlitchData0,
	      OutSignalName => "DATAOUT(0)",
	      OutTemp       => DATAOUT_zd(0),
	      Paths         => (
	      			0 => (CLOCK_ipd'last_event, tpd_CLOCK_DATAOUT_posedge(0), true),
				1 => (SLEEP_ipd'last_event, tpd_SLEEP_DATAOUT_posedge(0), true)
      			       ),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => DATAOUT(1),
	      GlitchData    => DATAOUT_GlitchData1,
	      OutSignalName => "DATAOUT(1)",
	      OutTemp       => DATAOUT_zd(1),
	      Paths         => (
	      			0 => (CLOCK_ipd'last_event, tpd_CLOCK_DATAOUT_posedge(1), true),
				1 => (SLEEP_ipd'last_event, tpd_SLEEP_DATAOUT_posedge(1), true)
      			       ),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => DATAOUT(2),
	      GlitchData    => DATAOUT_GlitchData2,
	      OutSignalName => "DATAOUT(2)",
	      OutTemp       => DATAOUT_zd(2),
	      Paths         => (
	      			0 => (CLOCK_ipd'last_event, tpd_CLOCK_DATAOUT_posedge(2), true),
				1 => (SLEEP_ipd'last_event, tpd_SLEEP_DATAOUT_posedge(2), true)
      			       ),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => DATAOUT(3),
	      GlitchData    => DATAOUT_GlitchData3,
	      OutSignalName => "DATAOUT(3)",
	      OutTemp       => DATAOUT_zd(3),
	      Paths         => (
	      			0 => (CLOCK_ipd'last_event, tpd_CLOCK_DATAOUT_posedge(3), true),
				1 => (SLEEP_ipd'last_event, tpd_SLEEP_DATAOUT_posedge(3), true)
      			       ),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => DATAOUT(4),
	      GlitchData    => DATAOUT_GlitchData4,
	      OutSignalName => "DATAOUT(4)",
	      OutTemp       => DATAOUT_zd(4),
	      Paths         => (
	      			0 => (CLOCK_ipd'last_event, tpd_CLOCK_DATAOUT_posedge(4), true),
				1 => (SLEEP_ipd'last_event, tpd_SLEEP_DATAOUT_posedge(4), true)
      			       ),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => DATAOUT(5),
	      GlitchData    => DATAOUT_GlitchData5,
	      OutSignalName => "DATAOUT(5)",
	      OutTemp       => DATAOUT_zd(5),
	      Paths         => (
	      			0 => (CLOCK_ipd'last_event, tpd_CLOCK_DATAOUT_posedge(5), true),
				1 => (SLEEP_ipd'last_event, tpd_SLEEP_DATAOUT_posedge(5), true)
      			       ),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => DATAOUT(6),
	      GlitchData    => DATAOUT_GlitchData6,
	      OutSignalName => "DATAOUT(6)",
	      OutTemp       => DATAOUT_zd(6),
	      Paths         => (
	      			0 => (CLOCK_ipd'last_event, tpd_CLOCK_DATAOUT_posedge(6), true),
				1 => (SLEEP_ipd'last_event, tpd_SLEEP_DATAOUT_posedge(6), true)
      			       ),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => DATAOUT(7),
	      GlitchData    => DATAOUT_GlitchData7,
	      OutSignalName => "DATAOUT(7)",
	      OutTemp       => DATAOUT_zd(7),
	      Paths         => (
	      			0 => (CLOCK_ipd'last_event, tpd_CLOCK_DATAOUT_posedge(7), true),
				1 => (SLEEP_ipd'last_event, tpd_SLEEP_DATAOUT_posedge(7), true)
      			       ),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => DATAOUT(8),
	      GlitchData    => DATAOUT_GlitchData8,
	      OutSignalName => "DATAOUT(8)",
	      OutTemp       => DATAOUT_zd(8),
	      Paths         => (
	      			0 => (CLOCK_ipd'last_event, tpd_CLOCK_DATAOUT_posedge(8), true),
				1 => (SLEEP_ipd'last_event, tpd_SLEEP_DATAOUT_posedge(8), true)
      			       ),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => DATAOUT(9),
	      GlitchData    => DATAOUT_GlitchData9,
	      OutSignalName => "DATAOUT(9)",
	      OutTemp       => DATAOUT_zd(9),
	      Paths         => (
	      			0 => (CLOCK_ipd'last_event, tpd_CLOCK_DATAOUT_posedge(9), true),
				1 => (SLEEP_ipd'last_event, tpd_SLEEP_DATAOUT_posedge(9), true)
      			       ),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => DATAOUT(10),
	      GlitchData    => DATAOUT_GlitchData10,
	      OutSignalName => "DATAOUT(10)",
	      OutTemp       => DATAOUT_zd(10),
	      Paths         => (
	      			0 => (CLOCK_ipd'last_event, tpd_CLOCK_DATAOUT_posedge(10), true),
				1 => (SLEEP_ipd'last_event, tpd_SLEEP_DATAOUT_posedge(10), true)
      			       ),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => DATAOUT(11),
	      GlitchData    => DATAOUT_GlitchData11,
	      OutSignalName => "DATAOUT(11)",
	      OutTemp       => DATAOUT_zd(11),
	      Paths         => (
	      			0 => (CLOCK_ipd'last_event, tpd_CLOCK_DATAOUT_posedge(11), true),
				1 => (SLEEP_ipd'last_event, tpd_SLEEP_DATAOUT_posedge(11), true)
      			       ),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => DATAOUT(12),
	      GlitchData    => DATAOUT_GlitchData12,
	      OutSignalName => "DATAOUT(12)",
	      OutTemp       => DATAOUT_zd(12),
	      Paths         => (
	      			0 => (CLOCK_ipd'last_event, tpd_CLOCK_DATAOUT_posedge(12), true),
				1 => (SLEEP_ipd'last_event, tpd_SLEEP_DATAOUT_posedge(12), true) ),
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => DATAOUT(13),
	      GlitchData    => DATAOUT_GlitchData13,
	      OutSignalName => "DATAOUT(13)",
	      OutTemp       => DATAOUT_zd(13),
	      Paths         => (
	      			0 => (CLOCK_ipd'last_event, tpd_CLOCK_DATAOUT_posedge(13), true),
				1 => (SLEEP_ipd'last_event, tpd_SLEEP_DATAOUT_posedge(13), true)
      			       ),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => DATAOUT(14),
	      GlitchData    => DATAOUT_GlitchData14,
	      OutSignalName => "DATAOUT(14)",
	      OutTemp       => DATAOUT_zd(14),
	      Paths         => (
	      			0 => (CLOCK_ipd'last_event, tpd_CLOCK_DATAOUT_posedge(14), true),
				1 => (SLEEP_ipd'last_event, tpd_SLEEP_DATAOUT_posedge(14), true)
      			       ),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	    VitalPathDelay01 (
	      OutSignal     => DATAOUT(15),
	      GlitchData    => DATAOUT_GlitchData15,
	      OutSignalName => "DATAOUT(15)",
	      OutTemp       => DATAOUT_zd(15),
	      Paths         => (
	      			0 => (CLOCK_ipd'last_event, tpd_CLOCK_DATAOUT_posedge(15), true),
				1 => (SLEEP_ipd'last_event, tpd_SLEEP_DATAOUT_posedge(15), true)
      			       ),
	      Mode          => OnEvent,
	      Xon           => Xon,
	      MsgOn         => MsgOn,
	      MsgSeverity   => warning);

	end process;

	end block;  	 
	
end SB_SPRAM256KA_V; 

------------------------------------------------------------------------
--					SB_IO_I3C
------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
--library	work;
use	work.std_logic_SBT.all;

entity	SB_IO_I3C is

	generic (
			NEG_TRIGGER : bit						:=	'0';
			PIN_TYPE	: bit_vector (5 downto 0)	:=	"000000";
			PULLUP		: bit						:=	'0';
			WEAK_PULLUP	: bit						:=  '0'; 
			IO_STANDARD	: string					:=	"SB_LVCMOS"
			);
	port 
		(
		D_OUT_1 		    : in std_logic;
		D_OUT_0 		    : in std_logic;
		CLOCK_ENABLE		: in std_logic;
		LATCH_INPUT_VALUE	: in std_logic;
		INPUT_CLK			: in std_logic;			
		D_IN_1				: out std_logic;
		D_IN_0				: out std_logic;
		OUTPUT_ENABLE		: in std_logic	:='H';
		OUTPUT_CLK			: in std_logic;			
		PU_ENB				: in std_logic ; 
		WEAK_PU_ENB			: in std_logic; 		
		PACKAGE_PIN			: inout	std_ulogic
		); 
		
end SB_IO_I3C ;

architecture SB_IO_I3C_V of SB_IO_I3C is

	component	preio_physical
	port	(
			hold	:	in 	std_logic;
			rstio	:	in	std_logic;
			bs_en	:	in	std_logic;
			shift	:	in	std_logic;
			tclk	:	in	std_logic;
			inclk	:	in	std_logic;
			outclk	:	in	std_logic;
			update	:	in	std_logic;
			oepin	:	in	std_logic;
			sdi		:	in	std_logic;
			mode	:	in	std_logic;
			hiz_b	:	in	std_logic;
			sdo		:	out	std_logic;
			dout1	:	out	std_logic;
			dout0	:	out	std_logic;
			ddr1	:	in	std_logic;
			ddr0	:	in	std_logic;
			padin	:	in	std_logic;
			padout	:	out	std_logic;
			padoen	:	out	std_logic;
			cbit	:	in	std_logic_vector	(5 downto 0)
			);
	end component;

	signal	inclk_n, outclk_n, inclk, outclk,sdo	:	std_logic;
	
	signal	bs_en	:	std_logic	:='0';	--Boundary scan enable           
	signal	shift	:	std_logic	:='0';	--Boundary scan shift            
	signal	tclk	:	std_logic	:='0';	--Boundary scan clock            
	signal	update	:	std_logic	:='0';	--Boundary scan update           
	signal	sdi		:	std_logic	:='0';	--Boundary scan serial data in   
	signal	mode	:	std_logic	:='0';	--Boundary scan mode             
	signal	hiz_b	:	std_logic	:='1';	--Boundary scan Tristate control 
	
	signal	pin_cbit:	std_logic_vector(5 downto 0);
	signal	neg_trig:	std_logic;
	signal	pull_up	:	std_logic;
	signal	hold,oepin,padoen,padout,padin	:	std_logic;
	signal INCLKE_sync , OUTCLKE_sync  	: std_logic;
	
	signal  net200 :	std_logic;
	
begin
	
	pin_cbit	<=	TO_STDLOGICVECTOR	(PIN_TYPE);
	neg_trig	<=	TO_STDLOGIC	(NEG_TRIGGER);
	pull_up		<=	TO_STDLOGIC	(PULLUP);

	inclk_n	<= 	INPUT_CLK xor neg_trig;
	outclk_n<=	OUTPUT_CLK xor neg_trig;
--	inclk	<=	inclk_n and CLOCK_ENABLE;
--	outclk	<=	outclk_n and CLOCK_ENABLE;

	net200 <= not(((not(PUENB) and PULLUP)  or ((not(WEAKPUENB) and WEAK_PULLUP))));
	
	process(inclk_n , CLOCK_ENABLE) is
         begin
                if(inclk_n ='0') then
                        INCLKE_sync  <= CLOCK_ENABLE;
                else
                        INCLKE_sync <= INCLKE_sync;
                end if ;
        end process;

        process(outclk_n , CLOCK_ENABLE) is
        begin
                if(outclk_n ='0') then
                        OUTCLKE_sync  <= CLOCK_ENABLE;
                else
                        OUTCLKE_sync <= OUTCLKE_sync;
                end if ;
        end process;

        inclk <= (inclk_n and INCLKE_sync);
        outclk <= (outclk_n and OUTCLKE_sync);
	
	hold	<=	LATCH_INPUT_VALUE;
	oepin	<=	OUTPUT_ENABLE;
	
	PACKAGE_PIN_i	:	process	(padoen, padout, PACKAGE_PIN)
	begin
		padin	<=	PACKAGE_PIN;
		if	(padoen='1') then
			PACKAGE_PIN	<=	'Z';
		else
			PACKAGE_PIN	<=	padout;
		end if;
	end process;
	
	PACKAGE_PIN_i_0:	process (net200, PACKAGE_PIN)
	begin
		if(net200='1') then
			PACKAGE_PIN <= 'Z';
		else 
			PACKAGE_PIN <= 'H';
		end if;
	end process;
	

-----------------------------------------------------------------	
	preio_physical_i	:	preio_physical
	port map	(
				hold	=>	hold,
				rstio	=>	'0',
				bs_en	=>	bs_en,
				shift	=>	shift,
				tclk	=>	tclk,
				inclk	=>	inclk,
				outclk	=>	outclk,
				update	=>	update,
				oepin	=>	oepin,
				sdi		=>	sdi,
				mode	=>	mode,
				hiz_b	=>	hiz_b,
				sdo		=>	sdo,
				dout1	=>	D_IN_1,
				dout0	=>	D_IN_0,
				ddr1	=>	D_OUT_1,
				ddr0	=>	D_OUT_0,
				padin	=>	padin,
				padout	=>	padout,
				padoen	=>	padoen,
				cbit	=>	pin_cbit
				);
end	SB_IO_I3C_V;

------------------------------------------------------------------------
--		SB_FILTER_50Ns 					     --
--  Glitch Filter with 50Ns Delay 				      -- 
------------------------------------------------------------------------


library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use IEEE.Vital_Primitives.all;
use IEEE.VITAL_Timing.all;

entity SB_FILTER_50NS is
  generic(
    Xon   : boolean := true;
    MsgOn : boolean := true;
   
      tipd_FILTERIN 		: VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_FILTERIN_FILTEROUT 	: VitalDelayType01 := (0.000 ns, 0.000 ns)
    );
  port(
    FILTEROUT : out std_logic;
    FILTERIN : in std_logic
    );
  attribute VITAL_LEVEL0 of SB_FILTER_50NS : entity is true;

end SB_FILTER_50NS;

architecture SB_FILTER_50NS_V  of SB_FILTER_50NS is
  attribute VITAL_LEVEL0 of SB_FILTER_50NS_V : architecture is true;

  signal FILTERIN_ipd : std_ulogic := 'X';
begin
  WireDelay : block
  begin
    VitalWireDelay (FILTERIN_ipd, FILTERIN, tipd_FILTERIN);
  end block;

  VITALBehavior           : process (FILTERIN_ipd)
    
      variable FILTEROUT_zd         : std_ulogic;
      variable FILTEROUT_GlitchData : VitalGlitchDataType;

    begin    

    FILTEROUT_zd := FILTERIN_ipd;


    VitalPathDelay01 (
      OutSignal     => FILTEROUT,
      GlitchData    => FILTEROUT_GlitchData,
      OutSignalName => "FILTEROUT",
      OutTemp       => FILTEROUT_zd,
      Paths         => (0 => (FILTERIN_ipd'last_event, tpd_FILTERIN_FILTEROUT, true)),
      Mode          => VitalTransport,
      Xon           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => warning);
  end process;
end SB_FILTER_50NS_V;






