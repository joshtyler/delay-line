// Top level module

module top(LED0, LED1);

output LED0, LED1;

//Hold LEDs
assign LED0 = 0;
assign LED1 = 1;

endmodule
